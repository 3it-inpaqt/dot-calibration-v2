* Netlist that describe the physical circuit (components and connexions between them) to simulate, in Xyce formalism.
* To make the translation from any network size, the circuit is scaled up automatically using Jinja template engine.
*
* Xyce: https://xyce.sandia.gov
* Jinja: https://jinja.palletsprojects.com

* ======================== Simulation parameters ==========================

.TRAN 0.30ns 331.00ns

* OPTIONS TIMEINT change the time integration parameters
* ERROPTION (If 0 Local Truncation Error is used)
* METHOD: Time integration method
* NLMIN, NLMAX:  lower and upper bound for the desired number of nonlinear iterations
* DELMAX: The maximum time step-size used
* This additional line allows to fix convergence problem but increases the simulation time
* List variables to save in the result table
.PRINT TRAN V(sum_h_out_003_001) V(hidden_activ_out_h003_001)
+ V(i_001) V(i_002) V(i_003) V(i_004) V(i_005) V(i_006) V(i_007) V(i_008) V(i_009) V(i_010) V(i_011) V(i_012) V(i_013) V(i_014) V(i_015) V(i_016) V(i_017) V(i_018) V(i_019) V(i_020) V(i_021) V(i_022) V(i_023) V(i_024) V(i_025) V(i_026) V(i_027) V(i_028) V(i_029) V(i_030) V(i_031) V(i_032) V(i_033) V(i_034) V(i_035) V(i_036) V(i_037) V(i_038) V(i_039) V(i_040) V(i_041) V(i_042) V(i_043) V(i_044) V(i_045) V(i_046) V(i_047) V(i_048) V(i_049) V(i_050) V(i_051) V(i_052) V(i_053) V(i_054) V(i_055) V(i_056) V(i_057) V(i_058) V(i_059) V(i_060) V(i_061) V(i_062) V(i_063) V(i_064)
+ V(sum_h_out_001_001) V(hidden_activ_out_h001_001) V(sum_h_out_001_002) V(hidden_activ_out_h001_002) V(sum_h_out_001_003) V(hidden_activ_out_h001_003) V(sum_h_out_001_004) V(hidden_activ_out_h001_004) V(sum_h_out_001_005) V(hidden_activ_out_h001_005) V(sum_h_out_001_006) V(hidden_activ_out_h001_006) V(sum_h_out_001_007) V(hidden_activ_out_h001_007) V(sum_h_out_001_008) V(hidden_activ_out_h001_008) V(sum_h_out_001_009) V(hidden_activ_out_h001_009) V(sum_h_out_001_010) V(hidden_activ_out_h001_010) V(sum_h_out_001_011) V(hidden_activ_out_h001_011) V(sum_h_out_001_012) V(hidden_activ_out_h001_012) V(sum_h_out_001_013) V(hidden_activ_out_h001_013) V(sum_h_out_001_014) V(hidden_activ_out_h001_014) V(sum_h_out_001_015) V(hidden_activ_out_h001_015) V(sum_h_out_001_016) V(hidden_activ_out_h001_016) V(sum_h_out_001_017) V(hidden_activ_out_h001_017) V(sum_h_out_001_018) V(hidden_activ_out_h001_018) V(sum_h_out_001_019) V(hidden_activ_out_h001_019) V(sum_h_out_001_020) V(hidden_activ_out_h001_020)
+ V(tia_h_out_001_001+) V(tia_h_out_001_001-) V(tia_h_out_001_002+) V(tia_h_out_001_002-) V(tia_h_out_001_003+) V(tia_h_out_001_003-) V(tia_h_out_001_004+) V(tia_h_out_001_004-) V(tia_h_out_001_005+) V(tia_h_out_001_005-) V(tia_h_out_001_006+) V(tia_h_out_001_006-) V(tia_h_out_001_007+) V(tia_h_out_001_007-) V(tia_h_out_001_008+) V(tia_h_out_001_008-) V(tia_h_out_001_009+) V(tia_h_out_001_009-) V(tia_h_out_001_010+) V(tia_h_out_001_010-) V(tia_h_out_001_011+) V(tia_h_out_001_011-) V(tia_h_out_001_012+) V(tia_h_out_001_012-) V(tia_h_out_001_013+) V(tia_h_out_001_013-) V(tia_h_out_001_014+) V(tia_h_out_001_014-) V(tia_h_out_001_015+) V(tia_h_out_001_015-) V(tia_h_out_001_016+) V(tia_h_out_001_016-) V(tia_h_out_001_017+) V(tia_h_out_001_017-) V(tia_h_out_001_018+) V(tia_h_out_001_018-) V(tia_h_out_001_019+) V(tia_h_out_001_019-) V(tia_h_out_001_020+) V(tia_h_out_001_020-)
+ V(b_001)
+ V(sum_h_out_002_001) V(hidden_activ_out_h002_001) V(sum_h_out_002_002) V(hidden_activ_out_h002_002) V(sum_h_out_002_003) V(hidden_activ_out_h002_003) V(sum_h_out_002_004) V(hidden_activ_out_h002_004) V(sum_h_out_002_005) V(hidden_activ_out_h002_005) V(sum_h_out_002_006) V(hidden_activ_out_h002_006) V(sum_h_out_002_007) V(hidden_activ_out_h002_007) V(sum_h_out_002_008) V(hidden_activ_out_h002_008) V(sum_h_out_002_009) V(hidden_activ_out_h002_009) V(sum_h_out_002_010) V(hidden_activ_out_h002_010)
+ V(tia_h_out_002_001+) V(tia_h_out_002_001-) V(tia_h_out_002_002+) V(tia_h_out_002_002-) V(tia_h_out_002_003+) V(tia_h_out_002_003-) V(tia_h_out_002_004+) V(tia_h_out_002_004-) V(tia_h_out_002_005+) V(tia_h_out_002_005-) V(tia_h_out_002_006+) V(tia_h_out_002_006-) V(tia_h_out_002_007+) V(tia_h_out_002_007-) V(tia_h_out_002_008+) V(tia_h_out_002_008-) V(tia_h_out_002_009+) V(tia_h_out_002_009-) V(tia_h_out_002_010+) V(tia_h_out_002_010-)
+ V(b_002)
+ V(sum_h_out_003_001) V(hidden_activ_out_h003_001)
+ V(tia_h_out_003_001+) V(tia_h_out_003_001-)
+ V(b_003)

* =============================== Models ==================================

* Call the defined components model from the specified path
*.INCLUDE "./components/MAX4223.sub"
.INCLUDE "./components/TLV3501.sub"
*.INCLUDE "./components/OPA684.sub"

* Import custom sub-circuits
.INCLUDE "./components/activations.sub"
.INCLUDE "./components/lumped_line.sub"
.INCLUDE "./components/Sigmoid3_HA.spice"

* Define diode model
.MODEL D_BAV74_1 D( IS=2.073F N=1 BV=50 IBV=100N RS=1.336 
+      CJO=2P VJ=750M M=330M FC=500M TT=5.771N 
+      EG=1.11 XTI=3 KF=0 AF=1 )

* ============================== Voltages =================================

* ----- Input pulses
* Vi_num: The input voltage as pulse sequences
Vi_001    i_001    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.083V 300.00ns 1.083V 301.00ns 0.950V
Vi_002    i_002    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.035V 300.00ns 1.035V 301.00ns 0.950V
Vi_003    i_003    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.000V 300.00ns 1.000V 301.00ns 0.950V
Vi_004    i_004    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.972V 300.00ns 0.972V 301.00ns 0.950V
Vi_005    i_005    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.009V 300.00ns 1.009V 301.00ns 0.950V
Vi_006    i_006    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.995V 300.00ns 0.995V 301.00ns 0.950V
Vi_007    i_007    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.042V 300.00ns 1.042V 301.00ns 0.950V
Vi_008    i_008    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.950V 300.00ns 0.950V 301.00ns 0.950V
Vi_009    i_009    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.080V 300.00ns 1.080V 301.00ns 0.950V
Vi_010    i_010    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.039V 300.00ns 1.039V 301.00ns 0.950V
Vi_011    i_011    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.995V 300.00ns 0.995V 301.00ns 0.950V
Vi_012    i_012    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.005V 300.00ns 1.005V 301.00ns 0.950V
Vi_013    i_013    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.010V 300.00ns 1.010V 301.00ns 0.950V
Vi_014    i_014    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.038V 300.00ns 1.038V 301.00ns 0.950V
Vi_015    i_015    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.053V 300.00ns 1.053V 301.00ns 0.950V
Vi_016    i_016    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.960V 300.00ns 0.960V 301.00ns 0.950V
Vi_017    i_017    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.073V 300.00ns 1.073V 301.00ns 0.950V
Vi_018    i_018    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.050V 300.00ns 1.050V 301.00ns 0.950V
Vi_019    i_019    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.992V 300.00ns 0.992V 301.00ns 0.950V
Vi_020    i_020    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.025V 300.00ns 1.025V 301.00ns 0.950V
Vi_021    i_021    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.072V 300.00ns 1.072V 301.00ns 0.950V
Vi_022    i_022    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.035V 300.00ns 1.035V 301.00ns 0.950V
Vi_023    i_023    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.081V 300.00ns 1.081V 301.00ns 0.950V
Vi_024    i_024    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.996V 300.00ns 0.996V 301.00ns 0.950V
Vi_025    i_025    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.104V 300.00ns 1.104V 301.00ns 0.950V
Vi_026    i_026    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.054V 300.00ns 1.054V 301.00ns 0.950V
Vi_027    i_027    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.019V 300.00ns 1.019V 301.00ns 0.950V
Vi_028    i_028    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.028V 300.00ns 1.028V 301.00ns 0.950V
Vi_029    i_029    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.034V 300.00ns 1.034V 301.00ns 0.950V
Vi_030    i_030    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.049V 300.00ns 1.049V 301.00ns 0.950V
Vi_031    i_031    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.072V 300.00ns 1.072V 301.00ns 0.950V
Vi_032    i_032    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.995V 300.00ns 0.995V 301.00ns 0.950V
Vi_033    i_033    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.130V 300.00ns 1.130V 301.00ns 0.950V
Vi_034    i_034    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.073V 300.00ns 1.073V 301.00ns 0.950V
Vi_035    i_035    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.030V 300.00ns 1.030V 301.00ns 0.950V
Vi_036    i_036    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.023V 300.00ns 1.023V 301.00ns 0.950V
Vi_037    i_037    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.087V 300.00ns 1.087V 301.00ns 0.950V
Vi_038    i_038    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.066V 300.00ns 1.066V 301.00ns 0.950V
Vi_039    i_039    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.086V 300.00ns 1.086V 301.00ns 0.950V
Vi_040    i_040    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.019V 300.00ns 1.019V 301.00ns 0.950V
Vi_041    i_041    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.150V 300.00ns 1.150V 301.00ns 0.950V
Vi_042    i_042    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.091V 300.00ns 1.091V 301.00ns 0.950V
Vi_043    i_043    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.036V 300.00ns 1.036V 301.00ns 0.950V
Vi_044    i_044    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.042V 300.00ns 1.042V 301.00ns 0.950V
Vi_045    i_045    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.094V 300.00ns 1.094V 301.00ns 0.950V
Vi_046    i_046    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.075V 300.00ns 1.075V 301.00ns 0.950V
Vi_047    i_047    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.103V 300.00ns 1.103V 301.00ns 0.950V
Vi_048    i_048    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.023V 300.00ns 1.023V 301.00ns 0.950V
Vi_049    i_049    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.136V 300.00ns 1.136V 301.00ns 0.950V
Vi_050    i_050    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.109V 300.00ns 1.109V 301.00ns 0.950V
Vi_051    i_051    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.062V 300.00ns 1.062V 301.00ns 0.950V
Vi_052    i_052    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.044V 300.00ns 1.044V 301.00ns 0.950V
Vi_053    i_053    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.100V 300.00ns 1.100V 301.00ns 0.950V
Vi_054    i_054    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.085V 300.00ns 1.085V 301.00ns 0.950V
Vi_055    i_055    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.091V 300.00ns 1.091V 301.00ns 0.950V
Vi_056    i_056    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.020V 300.00ns 1.020V 301.00ns 0.950V
Vi_057    i_057    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.133V 300.00ns 1.133V 301.00ns 0.950V
Vi_058    i_058    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.107V 300.00ns 1.107V 301.00ns 0.950V
Vi_059    i_059    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.074V 300.00ns 1.074V 301.00ns 0.950V
Vi_060    i_060    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.045V 300.00ns 1.045V 301.00ns 0.950V
Vi_061    i_061    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.115V 300.00ns 1.115V 301.00ns 0.950V
Vi_062    i_062    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.057V 300.00ns 1.057V 301.00ns 0.950V
Vi_063    i_063    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.135V 300.00ns 1.135V 301.00ns 0.950V
Vi_064    i_064    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.033V 300.00ns 1.033V 301.00ns 0.950V

* Vb_num: The bias voltage as pulse sequences

Vb_001    b_001    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.150V 300.00ns 1.150V 301.00ns 0.950V
Vb_002    b_002    0    PWL 0.00ns 0.950V 11.00ns 0.950V 12.00ns 1.150V 310.00ns 1.150V 311.00ns 0.950V
Vb_003    b_003    0    PWL 0.00ns 0.950V 21.00ns 0.950V 22.00ns 1.150V 320.00ns 1.150V 321.00ns 0.950V

Ve        Ve       0    3
Vcc-      Vcc-     0    -5
Vcc+      Vcc+     0    5

* ============================ NN Parameters ==============================
* Parameters (weights and bias) naming convention: "Rl_i_j+" where:
*   R: Always "R" to inform Xyce it is a resistance
*   l: layer name, "h" for the hidden and output layers and "b" for the biases.
*   i: index of the weight of a neuron (start from 1)
*   j: index of the neuron (start from 1)
*   +: parameter polarity, + or -

* ----------------------------- Layers -----------------------------


* ----- Weights
* Layer 001

* Neuron 1
Rh001_001_001+    i_001    tia_h_in_001_001+    121029.16352100707
Rh001_001_001-    i_001    tia_h_in_001_001-    26604.586298782495
Rh001_002_001+    i_002    tia_h_in_001_001+    120700.51264123355
Rh001_002_001-    i_002    tia_h_in_001_001-    23626.834583053416
Rh001_003_001+    i_003    tia_h_in_001_001+    99066.72376520271
Rh001_003_001-    i_003    tia_h_in_001_001-    118967.06792834178
Rh001_004_001+    i_004    tia_h_in_001_001+    27026.721587790697
Rh001_004_001-    i_004    tia_h_in_001_001-    120867.44497983945
Rh001_005_001+    i_005    tia_h_in_001_001+    23128.570645191023
Rh001_005_001-    i_005    tia_h_in_001_001-    120182.296121053
Rh001_006_001+    i_006    tia_h_in_001_001+    28828.173973941564
Rh001_006_001-    i_006    tia_h_in_001_001-    119932.69073462243
Rh001_007_001+    i_007    tia_h_in_001_001+    121200.46784558384
Rh001_007_001-    i_007    tia_h_in_001_001-    73781.3264762695
Rh001_008_001+    i_008    tia_h_in_001_001+    120934.83536510603
Rh001_008_001-    i_008    tia_h_in_001_001-    53878.36843904545
Rh001_009_001+    i_009    tia_h_in_001_001+    119915.71564731402
Rh001_009_001-    i_009    tia_h_in_001_001-    84535.00312183071
Rh001_010_001+    i_010    tia_h_in_001_001+    67166.7713389851
Rh001_010_001-    i_010    tia_h_in_001_001-    119800.99430376728
Rh001_011_001+    i_011    tia_h_in_001_001+    31113.384270098606
Rh001_011_001-    i_011    tia_h_in_001_001-    120557.91227530874
Rh001_012_001+    i_012    tia_h_in_001_001+    39248.35317571177
Rh001_012_001-    i_012    tia_h_in_001_001-    118378.32280535267
Rh001_013_001+    i_013    tia_h_in_001_001+    58584.1669905716
Rh001_013_001-    i_013    tia_h_in_001_001-    119015.94465609612
Rh001_014_001+    i_014    tia_h_in_001_001+    119597.50757370109
Rh001_014_001-    i_014    tia_h_in_001_001-    55363.16069077775
Rh001_015_001+    i_015    tia_h_in_001_001+    120107.8946401058
Rh001_015_001-    i_015    tia_h_in_001_001-    32021.3082161856
Rh001_016_001+    i_016    tia_h_in_001_001+    119293.88405307176
Rh001_016_001-    i_016    tia_h_in_001_001-    76841.54486013998
Rh001_017_001+    i_017    tia_h_in_001_001+    121210.730134822
Rh001_017_001-    i_017    tia_h_in_001_001-    55193.43296815773
Rh001_018_001+    i_018    tia_h_in_001_001+    42999.50704099807
Rh001_018_001-    i_018    tia_h_in_001_001-    119021.01688929688
Rh001_019_001+    i_019    tia_h_in_001_001+    5000
Rh001_019_001-    i_019    tia_h_in_001_001-    5000
Rh001_020_001+    i_020    tia_h_in_001_001+    27262.88979838742
Rh001_020_001-    i_020    tia_h_in_001_001-    121757.09400798022
Rh001_021_001+    i_021    tia_h_in_001_001+    88863.60024198492
Rh001_021_001-    i_021    tia_h_in_001_001-    118078.195521666
Rh001_022_001+    i_022    tia_h_in_001_001+    120597.82749383088
Rh001_022_001-    i_022    tia_h_in_001_001-    61897.82407518889
Rh001_023_001+    i_023    tia_h_in_001_001+    120321.632143572
Rh001_023_001-    i_023    tia_h_in_001_001-    66236.76090962837
Rh001_024_001+    i_024    tia_h_in_001_001+    5000
Rh001_024_001-    i_024    tia_h_in_001_001-    35429.4690051122
Rh001_025_001+    i_025    tia_h_in_001_001+    36682.87375241355
Rh001_025_001-    i_025    tia_h_in_001_001-    120620.47467524718
Rh001_026_001+    i_026    tia_h_in_001_001+    58177.69836784914
Rh001_026_001-    i_026    tia_h_in_001_001-    120016.38524913338
Rh001_027_001+    i_027    tia_h_in_001_001+    31207.98430624449
Rh001_027_001-    i_027    tia_h_in_001_001-    5000
Rh001_028_001+    i_028    tia_h_in_001_001+    94212.03532673832
Rh001_028_001-    i_028    tia_h_in_001_001-    121182.520665206
Rh001_029_001+    i_029    tia_h_in_001_001+    121167.23091797953
Rh001_029_001-    i_029    tia_h_in_001_001-    42080.19348379984
Rh001_030_001+    i_030    tia_h_in_001_001+    120755.44540835211
Rh001_030_001-    i_030    tia_h_in_001_001-    47473.507001308615
Rh001_031_001+    i_031    tia_h_in_001_001+    118991.45381286196
Rh001_031_001-    i_031    tia_h_in_001_001-    5000
Rh001_032_001+    i_032    tia_h_in_001_001+    70657.61542834865
Rh001_032_001-    i_032    tia_h_in_001_001-    121761.32525990887
Rh001_033_001+    i_033    tia_h_in_001_001+    5000
Rh001_033_001-    i_033    tia_h_in_001_001-    119201.21299929512
Rh001_034_001+    i_034    tia_h_in_001_001+    5000
Rh001_034_001-    i_034    tia_h_in_001_001-    117894.5906604111
Rh001_035_001+    i_035    tia_h_in_001_001+    119579.76800788291
Rh001_035_001-    i_035    tia_h_in_001_001-    111462.21723102785
Rh001_036_001+    i_036    tia_h_in_001_001+    119734.52330788861
Rh001_036_001-    i_036    tia_h_in_001_001-    91424.59199300379
Rh001_037_001+    i_037    tia_h_in_001_001+    119079.8457886117
Rh001_037_001-    i_037    tia_h_in_001_001-    81148.61874076909
Rh001_038_001+    i_038    tia_h_in_001_001+    121712.92325231015
Rh001_038_001-    i_038    tia_h_in_001_001-    5000
Rh001_039_001+    i_039    tia_h_in_001_001+    120724.87237827345
Rh001_039_001-    i_039    tia_h_in_001_001-    65864.45479272498
Rh001_040_001+    i_040    tia_h_in_001_001+    58519.2340798162
Rh001_040_001-    i_040    tia_h_in_001_001-    117883.57023549649
Rh001_041_001+    i_041    tia_h_in_001_001+    49104.64562337393
Rh001_041_001-    i_041    tia_h_in_001_001-    120404.56180774618
Rh001_042_001+    i_042    tia_h_in_001_001+    120819.15535247575
Rh001_042_001-    i_042    tia_h_in_001_001-    61352.60002885691
Rh001_043_001+    i_043    tia_h_in_001_001+    121084.919115528
Rh001_043_001-    i_043    tia_h_in_001_001-    114434.44467803476
Rh001_044_001+    i_044    tia_h_in_001_001+    120742.95807766056
Rh001_044_001-    i_044    tia_h_in_001_001-    120000
Rh001_045_001+    i_045    tia_h_in_001_001+    119715.57658638418
Rh001_045_001-    i_045    tia_h_in_001_001-    61786.62554168954
Rh001_046_001+    i_046    tia_h_in_001_001+    119401.62865622349
Rh001_046_001-    i_046    tia_h_in_001_001-    56250.88141116952
Rh001_047_001+    i_047    tia_h_in_001_001+    65559.40354338368
Rh001_047_001-    i_047    tia_h_in_001_001-    119387.64610584587
Rh001_048_001+    i_048    tia_h_in_001_001+    120000
Rh001_048_001-    i_048    tia_h_in_001_001-    121652.93046509744
Rh001_049_001+    i_049    tia_h_in_001_001+    46820.84422836565
Rh001_049_001-    i_049    tia_h_in_001_001-    120931.33951743871
Rh001_050_001+    i_050    tia_h_in_001_001+    45453.77177816445
Rh001_050_001-    i_050    tia_h_in_001_001-    120709.5452325173
Rh001_051_001+    i_051    tia_h_in_001_001+    120659.77217700976
Rh001_051_001-    i_051    tia_h_in_001_001-    88073.39375929406
Rh001_052_001+    i_052    tia_h_in_001_001+    120577.73638753795
Rh001_052_001-    i_052    tia_h_in_001_001-    57367.92204436632
Rh001_053_001+    i_053    tia_h_in_001_001+    119986.80195846618
Rh001_053_001-    i_053    tia_h_in_001_001-    43868.802307776175
Rh001_054_001+    i_054    tia_h_in_001_001+    121147.30264057912
Rh001_054_001-    i_054    tia_h_in_001_001-    5000
Rh001_055_001+    i_055    tia_h_in_001_001+    74914.91437249846
Rh001_055_001-    i_055    tia_h_in_001_001-    119963.17624841086
Rh001_056_001+    i_056    tia_h_in_001_001+    119229.75605637534
Rh001_056_001-    i_056    tia_h_in_001_001-    57366.91048877324
Rh001_057_001+    i_057    tia_h_in_001_001+    5000
Rh001_057_001-    i_057    tia_h_in_001_001-    120873.95309275421
Rh001_058_001+    i_058    tia_h_in_001_001+    120583.10870678225
Rh001_058_001-    i_058    tia_h_in_001_001-    84756.2913325527
Rh001_059_001+    i_059    tia_h_in_001_001+    121186.11766552611
Rh001_059_001-    i_059    tia_h_in_001_001-    21599.157981302662
Rh001_060_001+    i_060    tia_h_in_001_001+    120000
Rh001_060_001-    i_060    tia_h_in_001_001-    22381.546298514422
Rh001_061_001+    i_061    tia_h_in_001_001+    120528.75078643013
Rh001_061_001-    i_061    tia_h_in_001_001-    101128.58965972858
Rh001_062_001+    i_062    tia_h_in_001_001+    40198.465110336445
Rh001_062_001-    i_062    tia_h_in_001_001-    122257.77731796815
Rh001_063_001+    i_063    tia_h_in_001_001+    27886.41399205122
Rh001_063_001-    i_063    tia_h_in_001_001-    120469.91563692568
Rh001_064_001+    i_064    tia_h_in_001_001+    33078.534065266096
Rh001_064_001-    i_064    tia_h_in_001_001-    119897.59028799438

* Neuron 2
Rh001_001_002+    i_001    tia_h_in_001_002+    120118.86553775534
Rh001_001_002-    i_001    tia_h_in_001_002-    31893.397836213906
Rh001_002_002+    i_002    tia_h_in_001_002+    119930.54450732902
Rh001_002_002-    i_002    tia_h_in_001_002-    28570.73519517037
Rh001_003_002+    i_003    tia_h_in_001_002+    119901.97769094586
Rh001_003_002-    i_003    tia_h_in_001_002-    55736.077821823266
Rh001_004_002+    i_004    tia_h_in_001_002+    121302.1012975004
Rh001_004_002-    i_004    tia_h_in_001_002-    5000
Rh001_005_002+    i_005    tia_h_in_001_002+    117596.08690476384
Rh001_005_002-    i_005    tia_h_in_001_002-    63596.146984324085
Rh001_006_002+    i_006    tia_h_in_001_002+    118908.30794247072
Rh001_006_002-    i_006    tia_h_in_001_002-    33179.966503976
Rh001_007_002+    i_007    tia_h_in_001_002+    120182.18356661846
Rh001_007_002-    i_007    tia_h_in_001_002-    29716.475908658893
Rh001_008_002+    i_008    tia_h_in_001_002+    120147.01246091303
Rh001_008_002-    i_008    tia_h_in_001_002-    35151.18518860717
Rh001_009_002+    i_009    tia_h_in_001_002+    121343.47366748034
Rh001_009_002-    i_009    tia_h_in_001_002-    26188.032196971817
Rh001_010_002+    i_010    tia_h_in_001_002+    43237.330392619464
Rh001_010_002-    i_010    tia_h_in_001_002-    120000
Rh001_011_002+    i_011    tia_h_in_001_002+    119826.64171868587
Rh001_011_002-    i_011    tia_h_in_001_002-    75404.42100094547
Rh001_012_002+    i_012    tia_h_in_001_002+    41256.94270631952
Rh001_012_002-    i_012    tia_h_in_001_002-    121670.88667425285
Rh001_013_002+    i_013    tia_h_in_001_002+    99340.10547055124
Rh001_013_002-    i_013    tia_h_in_001_002-    120467.52955585823
Rh001_014_002+    i_014    tia_h_in_001_002+    119243.11334466447
Rh001_014_002-    i_014    tia_h_in_001_002-    101298.81485079302
Rh001_015_002+    i_015    tia_h_in_001_002+    56601.57084304448
Rh001_015_002-    i_015    tia_h_in_001_002-    119009.83536056962
Rh001_016_002+    i_016    tia_h_in_001_002+    63458.81162971003
Rh001_016_002-    i_016    tia_h_in_001_002-    120590.1559381146
Rh001_017_002+    i_017    tia_h_in_001_002+    30750.904686822712
Rh001_017_002-    i_017    tia_h_in_001_002-    121024.19092412459
Rh001_018_002+    i_018    tia_h_in_001_002+    118835.99910084043
Rh001_018_002-    i_018    tia_h_in_001_002-    5000
Rh001_019_002+    i_019    tia_h_in_001_002+    113449.80559516042
Rh001_019_002-    i_019    tia_h_in_001_002-    119897.81702165559
Rh001_020_002+    i_020    tia_h_in_001_002+    119584.87828560824
Rh001_020_002-    i_020    tia_h_in_001_002-    66826.95548673034
Rh001_021_002+    i_021    tia_h_in_001_002+    87508.82974697194
Rh001_021_002-    i_021    tia_h_in_001_002-    5000
Rh001_022_002+    i_022    tia_h_in_001_002+    37846.835835416096
Rh001_022_002-    i_022    tia_h_in_001_002-    119904.43629330829
Rh001_023_002+    i_023    tia_h_in_001_002+    27537.280127937134
Rh001_023_002-    i_023    tia_h_in_001_002-    119876.68191365177
Rh001_024_002+    i_024    tia_h_in_001_002+    25895.043599129433
Rh001_024_002-    i_024    tia_h_in_001_002-    120431.42344625675
Rh001_025_002+    i_025    tia_h_in_001_002+    53400.127319347885
Rh001_025_002-    i_025    tia_h_in_001_002-    5000
Rh001_026_002+    i_026    tia_h_in_001_002+    51519.2361083474
Rh001_026_002-    i_026    tia_h_in_001_002-    121506.54590763112
Rh001_027_002+    i_027    tia_h_in_001_002+    120762.31704315446
Rh001_027_002-    i_027    tia_h_in_001_002-    58256.769572446945
Rh001_028_002+    i_028    tia_h_in_001_002+    120960.13649939174
Rh001_028_002-    i_028    tia_h_in_001_002-    51488.761166624245
Rh001_029_002+    i_029    tia_h_in_001_002+    37841.995390097174
Rh001_029_002-    i_029    tia_h_in_001_002-    120930.71608948539
Rh001_030_002+    i_030    tia_h_in_001_002+    78557.22596637617
Rh001_030_002-    i_030    tia_h_in_001_002-    121919.91858830338
Rh001_031_002+    i_031    tia_h_in_001_002+    86243.34497664182
Rh001_031_002-    i_031    tia_h_in_001_002-    121372.53772876457
Rh001_032_002+    i_032    tia_h_in_001_002+    117629.28786533677
Rh001_032_002-    i_032    tia_h_in_001_002-    118978.59967686764
Rh001_033_002+    i_033    tia_h_in_001_002+    5000
Rh001_033_002-    i_033    tia_h_in_001_002-    119337.56261455132
Rh001_034_002+    i_034    tia_h_in_001_002+    55371.334880438895
Rh001_034_002-    i_034    tia_h_in_001_002-    5000
Rh001_035_002+    i_035    tia_h_in_001_002+    94669.56005628883
Rh001_035_002-    i_035    tia_h_in_001_002-    120284.07619211814
Rh001_036_002+    i_036    tia_h_in_001_002+    119779.26400485195
Rh001_036_002-    i_036    tia_h_in_001_002-    80534.49958293657
Rh001_037_002+    i_037    tia_h_in_001_002+    95082.5894970481
Rh001_037_002-    i_037    tia_h_in_001_002-    119507.93851797601
Rh001_038_002+    i_038    tia_h_in_001_002+    120163.810515824
Rh001_038_002-    i_038    tia_h_in_001_002-    70799.91047134368
Rh001_039_002+    i_039    tia_h_in_001_002+    120000
Rh001_039_002-    i_039    tia_h_in_001_002-    36830.27157437423
Rh001_040_002+    i_040    tia_h_in_001_002+    119360.86493603843
Rh001_040_002-    i_040    tia_h_in_001_002-    54575.51638461993
Rh001_041_002+    i_041    tia_h_in_001_002+    102522.56601684052
Rh001_041_002-    i_041    tia_h_in_001_002-    119552.94720866633
Rh001_042_002+    i_042    tia_h_in_001_002+    59608.534336693505
Rh001_042_002-    i_042    tia_h_in_001_002-    119447.60364910704
Rh001_043_002+    i_043    tia_h_in_001_002+    33263.64300092399
Rh001_043_002-    i_043    tia_h_in_001_002-    118693.33637250277
Rh001_044_002+    i_044    tia_h_in_001_002+    54201.70566578236
Rh001_044_002-    i_044    tia_h_in_001_002-    119956.40352209842
Rh001_045_002+    i_045    tia_h_in_001_002+    122836.19026190935
Rh001_045_002-    i_045    tia_h_in_001_002-    40600.337870123185
Rh001_046_002+    i_046    tia_h_in_001_002+    120701.52665218673
Rh001_046_002-    i_046    tia_h_in_001_002-    37884.659014952
Rh001_047_002+    i_047    tia_h_in_001_002+    120755.21380744262
Rh001_047_002-    i_047    tia_h_in_001_002-    71995.58251576943
Rh001_048_002+    i_048    tia_h_in_001_002+    120673.35468967493
Rh001_048_002-    i_048    tia_h_in_001_002-    82195.36838234804
Rh001_049_002+    i_049    tia_h_in_001_002+    118669.65498598573
Rh001_049_002-    i_049    tia_h_in_001_002-    50561.3833940703
Rh001_050_002+    i_050    tia_h_in_001_002+    117926.27405934242
Rh001_050_002-    i_050    tia_h_in_001_002-    92553.31410539684
Rh001_051_002+    i_051    tia_h_in_001_002+    118776.43971685552
Rh001_051_002-    i_051    tia_h_in_001_002-    82146.95683906639
Rh001_052_002+    i_052    tia_h_in_001_002+    120064.14512474021
Rh001_052_002-    i_052    tia_h_in_001_002-    91403.23958384457
Rh001_053_002+    i_053    tia_h_in_001_002+    121523.25805450027
Rh001_053_002-    i_053    tia_h_in_001_002-    80429.58020959025
Rh001_054_002+    i_054    tia_h_in_001_002+    54172.146330492236
Rh001_054_002-    i_054    tia_h_in_001_002-    119270.79835197376
Rh001_055_002+    i_055    tia_h_in_001_002+    120000
Rh001_055_002-    i_055    tia_h_in_001_002-    61229.19126031693
Rh001_056_002+    i_056    tia_h_in_001_002+    120577.35462419187
Rh001_056_002-    i_056    tia_h_in_001_002-    120000
Rh001_057_002+    i_057    tia_h_in_001_002+    122052.60758120246
Rh001_057_002-    i_057    tia_h_in_001_002-    5000
Rh001_058_002+    i_058    tia_h_in_001_002+    121098.95493620756
Rh001_058_002-    i_058    tia_h_in_001_002-    98693.05793021836
Rh001_059_002+    i_059    tia_h_in_001_002+    120257.75305601688
Rh001_059_002-    i_059    tia_h_in_001_002-    57253.80707325487
Rh001_060_002+    i_060    tia_h_in_001_002+    120969.00855613276
Rh001_060_002-    i_060    tia_h_in_001_002-    108728.48898013277
Rh001_061_002+    i_061    tia_h_in_001_002+    120000
Rh001_061_002-    i_061    tia_h_in_001_002-    119837.39796414689
Rh001_062_002+    i_062    tia_h_in_001_002+    72816.68134412458
Rh001_062_002-    i_062    tia_h_in_001_002-    119423.60623205609
Rh001_063_002+    i_063    tia_h_in_001_002+    5000
Rh001_063_002-    i_063    tia_h_in_001_002-    119446.52748243276
Rh001_064_002+    i_064    tia_h_in_001_002+    119073.58972069657
Rh001_064_002-    i_064    tia_h_in_001_002-    56740.36826677557

* Neuron 3
Rh001_001_003+    i_001    tia_h_in_001_003+    121281.7900333057
Rh001_001_003-    i_001    tia_h_in_001_003-    53868.30956484281
Rh001_002_003+    i_002    tia_h_in_001_003+    120845.06337933675
Rh001_002_003-    i_002    tia_h_in_001_003-    62371.400567458666
Rh001_003_003+    i_003    tia_h_in_001_003+    28030.444210011054
Rh001_003_003-    i_003    tia_h_in_001_003-    119897.91445131891
Rh001_004_003+    i_004    tia_h_in_001_003+    18105.73496034543
Rh001_004_003-    i_004    tia_h_in_001_003-    120805.06827609563
Rh001_005_003+    i_005    tia_h_in_001_003+    35792.48693603936
Rh001_005_003-    i_005    tia_h_in_001_003-    120148.55147328491
Rh001_006_003+    i_006    tia_h_in_001_003+    118210.94046188564
Rh001_006_003-    i_006    tia_h_in_001_003-    81928.80438374521
Rh001_007_003+    i_007    tia_h_in_001_003+    120331.87516238283
Rh001_007_003-    i_007    tia_h_in_001_003-    43823.62860770307
Rh001_008_003+    i_008    tia_h_in_001_003+    120000
Rh001_008_003-    i_008    tia_h_in_001_003-    21518.756767480856
Rh001_009_003+    i_009    tia_h_in_001_003+    120000
Rh001_009_003-    i_009    tia_h_in_001_003-    119240.42074844263
Rh001_010_003+    i_010    tia_h_in_001_003+    49170.10553222382
Rh001_010_003-    i_010    tia_h_in_001_003-    121173.10020593874
Rh001_011_003+    i_011    tia_h_in_001_003+    41106.76903689421
Rh001_011_003-    i_011    tia_h_in_001_003-    120088.05141155767
Rh001_012_003+    i_012    tia_h_in_001_003+    121139.47070562915
Rh001_012_003-    i_012    tia_h_in_001_003-    71404.26913499692
Rh001_013_003+    i_013    tia_h_in_001_003+    5000
Rh001_013_003-    i_013    tia_h_in_001_003-    105545.56891823615
Rh001_014_003+    i_014    tia_h_in_001_003+    118592.77171113857
Rh001_014_003-    i_014    tia_h_in_001_003-    50674.76528979615
Rh001_015_003+    i_015    tia_h_in_001_003+    118455.13614281775
Rh001_015_003-    i_015    tia_h_in_001_003-    45042.478193923955
Rh001_016_003+    i_016    tia_h_in_001_003+    119568.01474934634
Rh001_016_003-    i_016    tia_h_in_001_003-    74299.74505447646
Rh001_017_003+    i_017    tia_h_in_001_003+    69454.59596904038
Rh001_017_003-    i_017    tia_h_in_001_003-    120553.73592553234
Rh001_018_003+    i_018    tia_h_in_001_003+    60781.59575496167
Rh001_018_003-    i_018    tia_h_in_001_003-    119985.87957207485
Rh001_019_003+    i_019    tia_h_in_001_003+    32928.269136970695
Rh001_019_003-    i_019    tia_h_in_001_003-    120855.14847580975
Rh001_020_003+    i_020    tia_h_in_001_003+    75040.06885422367
Rh001_020_003-    i_020    tia_h_in_001_003-    121236.19420223539
Rh001_021_003+    i_021    tia_h_in_001_003+    117743.85500516628
Rh001_021_003-    i_021    tia_h_in_001_003-    120039.83387006266
Rh001_022_003+    i_022    tia_h_in_001_003+    120448.32912951487
Rh001_022_003-    i_022    tia_h_in_001_003-    43580.345693074705
Rh001_023_003+    i_023    tia_h_in_001_003+    121968.1851077348
Rh001_023_003-    i_023    tia_h_in_001_003-    54073.38655183732
Rh001_024_003+    i_024    tia_h_in_001_003+    118239.06543487968
Rh001_024_003-    i_024    tia_h_in_001_003-    55360.91161302506
Rh001_025_003+    i_025    tia_h_in_001_003+    38660.395074076434
Rh001_025_003-    i_025    tia_h_in_001_003-    119734.3468821704
Rh001_026_003+    i_026    tia_h_in_001_003+    58100.9187858976
Rh001_026_003-    i_026    tia_h_in_001_003-    120197.0691992553
Rh001_027_003+    i_027    tia_h_in_001_003+    74610.55370243029
Rh001_027_003-    i_027    tia_h_in_001_003-    121504.66331986028
Rh001_028_003+    i_028    tia_h_in_001_003+    119775.92880606535
Rh001_028_003-    i_028    tia_h_in_001_003-    42197.68594932652
Rh001_029_003+    i_029    tia_h_in_001_003+    120035.23166915501
Rh001_029_003-    i_029    tia_h_in_001_003-    72446.59187047115
Rh001_030_003+    i_030    tia_h_in_001_003+    119620.72226204941
Rh001_030_003-    i_030    tia_h_in_001_003-    71344.8496475117
Rh001_031_003+    i_031    tia_h_in_001_003+    81751.11077804567
Rh001_031_003-    i_031    tia_h_in_001_003-    120921.236606053
Rh001_032_003+    i_032    tia_h_in_001_003+    71533.93587646786
Rh001_032_003-    i_032    tia_h_in_001_003-    118706.20844748613
Rh001_033_003+    i_033    tia_h_in_001_003+    55495.84697926304
Rh001_033_003-    i_033    tia_h_in_001_003-    119897.62023254871
Rh001_034_003+    i_034    tia_h_in_001_003+    120000
Rh001_034_003-    i_034    tia_h_in_001_003-    118445.983627359
Rh001_035_003+    i_035    tia_h_in_001_003+    119892.57407670822
Rh001_035_003-    i_035    tia_h_in_001_003-    42612.46503199381
Rh001_036_003+    i_036    tia_h_in_001_003+    5000
Rh001_036_003-    i_036    tia_h_in_001_003-    62293.398674073476
Rh001_037_003+    i_037    tia_h_in_001_003+    120810.12247335582
Rh001_037_003-    i_037    tia_h_in_001_003-    87984.50372526102
Rh001_038_003+    i_038    tia_h_in_001_003+    120699.3275160681
Rh001_038_003-    i_038    tia_h_in_001_003-    55519.599407762034
Rh001_039_003+    i_039    tia_h_in_001_003+    93375.15399101653
Rh001_039_003-    i_039    tia_h_in_001_003-    121027.68060512267
Rh001_040_003+    i_040    tia_h_in_001_003+    33281.79673825481
Rh001_040_003-    i_040    tia_h_in_001_003-    120431.24831279856
Rh001_041_003+    i_041    tia_h_in_001_003+    80159.88340668194
Rh001_041_003-    i_041    tia_h_in_001_003-    120909.77889840507
Rh001_042_003+    i_042    tia_h_in_001_003+    119380.73304435522
Rh001_042_003-    i_042    tia_h_in_001_003-    109446.95375581965
Rh001_043_003+    i_043    tia_h_in_001_003+    119389.95619458554
Rh001_043_003-    i_043    tia_h_in_001_003-    46168.03502808197
Rh001_044_003+    i_044    tia_h_in_001_003+    119605.74262362554
Rh001_044_003-    i_044    tia_h_in_001_003-    75505.19752374223
Rh001_045_003+    i_045    tia_h_in_001_003+    119494.4988313774
Rh001_045_003-    i_045    tia_h_in_001_003-    76611.29653142496
Rh001_046_003+    i_046    tia_h_in_001_003+    91777.87865734682
Rh001_046_003-    i_046    tia_h_in_001_003-    120594.54926445114
Rh001_047_003+    i_047    tia_h_in_001_003+    31252.99633975177
Rh001_047_003-    i_047    tia_h_in_001_003-    120704.76753851162
Rh001_048_003+    i_048    tia_h_in_001_003+    33459.0817827607
Rh001_048_003-    i_048    tia_h_in_001_003-    120824.07221878743
Rh001_049_003+    i_049    tia_h_in_001_003+    77449.55264341984
Rh001_049_003-    i_049    tia_h_in_001_003-    120232.45001087985
Rh001_050_003+    i_050    tia_h_in_001_003+    118219.43535663912
Rh001_050_003-    i_050    tia_h_in_001_003-    120000
Rh001_051_003+    i_051    tia_h_in_001_003+    118458.01052511386
Rh001_051_003-    i_051    tia_h_in_001_003-    91678.06542479954
Rh001_052_003+    i_052    tia_h_in_001_003+    118918.18864451058
Rh001_052_003-    i_052    tia_h_in_001_003-    58743.65080166038
Rh001_053_003+    i_053    tia_h_in_001_003+    120089.93170545784
Rh001_053_003-    i_053    tia_h_in_001_003-    44650.87213520809
Rh001_054_003+    i_054    tia_h_in_001_003+    121450.0034254852
Rh001_054_003-    i_054    tia_h_in_001_003-    70572.86561137455
Rh001_055_003+    i_055    tia_h_in_001_003+    40021.31541510039
Rh001_055_003-    i_055    tia_h_in_001_003-    121492.83629782023
Rh001_056_003+    i_056    tia_h_in_001_003+    72173.4309089441
Rh001_056_003-    i_056    tia_h_in_001_003-    120256.07237554081
Rh001_057_003+    i_057    tia_h_in_001_003+    120868.43143363748
Rh001_057_003-    i_057    tia_h_in_001_003-    35218.64132279253
Rh001_058_003+    i_058    tia_h_in_001_003+    120627.25824202002
Rh001_058_003-    i_058    tia_h_in_001_003-    47351.756769717176
Rh001_059_003+    i_059    tia_h_in_001_003+    120000
Rh001_059_003-    i_059    tia_h_in_001_003-    31731.489127195204
Rh001_060_003+    i_060    tia_h_in_001_003+    121570.39241875554
Rh001_060_003-    i_060    tia_h_in_001_003-    120000
Rh001_061_003+    i_061    tia_h_in_001_003+    49960.72412366511
Rh001_061_003-    i_061    tia_h_in_001_003-    5000
Rh001_062_003+    i_062    tia_h_in_001_003+    19931.964763492433
Rh001_062_003-    i_062    tia_h_in_001_003-    120601.80831275754
Rh001_063_003+    i_063    tia_h_in_001_003+    49294.309378572056
Rh001_063_003-    i_063    tia_h_in_001_003-    119370.57171931448
Rh001_064_003+    i_064    tia_h_in_001_003+    68783.56388801732
Rh001_064_003-    i_064    tia_h_in_001_003-    120427.08988300283

* Neuron 4
Rh001_001_004+    i_001    tia_h_in_001_004+    118584.68690874074
Rh001_001_004-    i_001    tia_h_in_001_004-    5000
Rh001_002_004+    i_002    tia_h_in_001_004+    120541.03434549714
Rh001_002_004-    i_002    tia_h_in_001_004-    102903.8005075605
Rh001_003_004+    i_003    tia_h_in_001_004+    5000
Rh001_003_004-    i_003    tia_h_in_001_004-    119202.11645986706
Rh001_004_004+    i_004    tia_h_in_001_004+    93701.5336439877
Rh001_004_004-    i_004    tia_h_in_001_004-    119660.75128075885
Rh001_005_004+    i_005    tia_h_in_001_004+    119454.22933784332
Rh001_005_004-    i_005    tia_h_in_001_004-    53817.77876801831
Rh001_006_004+    i_006    tia_h_in_001_004+    118900.94706945562
Rh001_006_004-    i_006    tia_h_in_001_004-    78340.9900399082
Rh001_007_004+    i_007    tia_h_in_001_004+    60488.841980498524
Rh001_007_004-    i_007    tia_h_in_001_004-    121138.64984182794
Rh001_008_004+    i_008    tia_h_in_001_004+    86361.25044661909
Rh001_008_004-    i_008    tia_h_in_001_004-    118453.60050897753
Rh001_009_004+    i_009    tia_h_in_001_004+    119577.80772915934
Rh001_009_004-    i_009    tia_h_in_001_004-    105600.94672379477
Rh001_010_004+    i_010    tia_h_in_001_004+    118691.80233023832
Rh001_010_004-    i_010    tia_h_in_001_004-    64647.94599115415
Rh001_011_004+    i_011    tia_h_in_001_004+    120775.38960135299
Rh001_011_004-    i_011    tia_h_in_001_004-    65018.999287999504
Rh001_012_004+    i_012    tia_h_in_001_004+    119961.97416760527
Rh001_012_004-    i_012    tia_h_in_001_004-    55089.62134170359
Rh001_013_004+    i_013    tia_h_in_001_004+    119761.75731152252
Rh001_013_004-    i_013    tia_h_in_001_004-    80869.17621083882
Rh001_014_004+    i_014    tia_h_in_001_004+    90073.6137952175
Rh001_014_004-    i_014    tia_h_in_001_004-    118612.14996019876
Rh001_015_004+    i_015    tia_h_in_001_004+    70430.26785764712
Rh001_015_004-    i_015    tia_h_in_001_004-    119114.81576574322
Rh001_016_004+    i_016    tia_h_in_001_004+    81310.69654073598
Rh001_016_004-    i_016    tia_h_in_001_004-    118623.21364922052
Rh001_017_004+    i_017    tia_h_in_001_004+    121693.1256258482
Rh001_017_004-    i_017    tia_h_in_001_004-    54519.45691934599
Rh001_018_004+    i_018    tia_h_in_001_004+    120318.18791974221
Rh001_018_004-    i_018    tia_h_in_001_004-    65094.62886888628
Rh001_019_004+    i_019    tia_h_in_001_004+    119157.08143921403
Rh001_019_004-    i_019    tia_h_in_001_004-    5000
Rh001_020_004+    i_020    tia_h_in_001_004+    55895.88952922315
Rh001_020_004-    i_020    tia_h_in_001_004-    120000
Rh001_021_004+    i_021    tia_h_in_001_004+    108437.1758381001
Rh001_021_004-    i_021    tia_h_in_001_004-    119834.73880236523
Rh001_022_004+    i_022    tia_h_in_001_004+    119872.4223474908
Rh001_022_004-    i_022    tia_h_in_001_004-    83398.50505622727
Rh001_023_004+    i_023    tia_h_in_001_004+    83943.71123929799
Rh001_023_004-    i_023    tia_h_in_001_004-    119972.92873064804
Rh001_024_004+    i_024    tia_h_in_001_004+    119791.88078068038
Rh001_024_004-    i_024    tia_h_in_001_004-    75279.50658495341
Rh001_025_004+    i_025    tia_h_in_001_004+    119370.66736284165
Rh001_025_004-    i_025    tia_h_in_001_004-    62912.221178478685
Rh001_026_004+    i_026    tia_h_in_001_004+    65087.49598155228
Rh001_026_004-    i_026    tia_h_in_001_004-    119484.61965595538
Rh001_027_004+    i_027    tia_h_in_001_004+    119207.85828433344
Rh001_027_004-    i_027    tia_h_in_001_004-    73013.89482699535
Rh001_028_004+    i_028    tia_h_in_001_004+    121178.48764683922
Rh001_028_004-    i_028    tia_h_in_001_004-    90478.34214022841
Rh001_029_004+    i_029    tia_h_in_001_004+    119062.77571562918
Rh001_029_004-    i_029    tia_h_in_001_004-    51583.155379144475
Rh001_030_004+    i_030    tia_h_in_001_004+    5000
Rh001_030_004-    i_030    tia_h_in_001_004-    119685.01028299969
Rh001_031_004+    i_031    tia_h_in_001_004+    64603.21365391724
Rh001_031_004-    i_031    tia_h_in_001_004-    121559.84031608904
Rh001_032_004+    i_032    tia_h_in_001_004+    87312.84656208965
Rh001_032_004-    i_032    tia_h_in_001_004-    119613.80750527783
Rh001_033_004+    i_033    tia_h_in_001_004+    120224.35460059273
Rh001_033_004-    i_033    tia_h_in_001_004-    60924.738448159405
Rh001_034_004+    i_034    tia_h_in_001_004+    120162.13541787698
Rh001_034_004-    i_034    tia_h_in_001_004-    51605.03682516693
Rh001_035_004+    i_035    tia_h_in_001_004+    119258.59065701236
Rh001_035_004-    i_035    tia_h_in_001_004-    58130.98237283838
Rh001_036_004+    i_036    tia_h_in_001_004+    65388.907583762826
Rh001_036_004-    i_036    tia_h_in_001_004-    121699.81087114614
Rh001_037_004+    i_037    tia_h_in_001_004+    5000
Rh001_037_004-    i_037    tia_h_in_001_004-    117895.14963400425
Rh001_038_004+    i_038    tia_h_in_001_004+    60504.99252983953
Rh001_038_004-    i_038    tia_h_in_001_004-    119374.15604075725
Rh001_039_004+    i_039    tia_h_in_001_004+    120000
Rh001_039_004-    i_039    tia_h_in_001_004-    119872.93054640335
Rh001_040_004+    i_040    tia_h_in_001_004+    98823.06992346016
Rh001_040_004-    i_040    tia_h_in_001_004-    120486.67601782865
Rh001_041_004+    i_041    tia_h_in_001_004+    119590.4749670415
Rh001_041_004-    i_041    tia_h_in_001_004-    109752.41953901234
Rh001_042_004+    i_042    tia_h_in_001_004+    119700.72538248694
Rh001_042_004-    i_042    tia_h_in_001_004-    59024.103684094494
Rh001_043_004+    i_043    tia_h_in_001_004+    121085.36781020906
Rh001_043_004-    i_043    tia_h_in_001_004-    56414.41882760754
Rh001_044_004+    i_044    tia_h_in_001_004+    120235.46661536915
Rh001_044_004-    i_044    tia_h_in_001_004-    54021.817093250975
Rh001_045_004+    i_045    tia_h_in_001_004+    81871.08921111713
Rh001_045_004-    i_045    tia_h_in_001_004-    120997.99071642355
Rh001_046_004+    i_046    tia_h_in_001_004+    120814.92199982813
Rh001_046_004-    i_046    tia_h_in_001_004-    70585.992552786
Rh001_047_004+    i_047    tia_h_in_001_004+    120790.12658533169
Rh001_047_004-    i_047    tia_h_in_001_004-    89534.58868168997
Rh001_048_004+    i_048    tia_h_in_001_004+    120000
Rh001_048_004-    i_048    tia_h_in_001_004-    66590.61640393037
Rh001_049_004+    i_049    tia_h_in_001_004+    119061.08163771093
Rh001_049_004-    i_049    tia_h_in_001_004-    90073.92290065545
Rh001_050_004+    i_050    tia_h_in_001_004+    120097.87984150174
Rh001_050_004-    i_050    tia_h_in_001_004-    61136.926535750004
Rh001_051_004+    i_051    tia_h_in_001_004+    119260.43164470559
Rh001_051_004-    i_051    tia_h_in_001_004-    63899.49713488776
Rh001_052_004+    i_052    tia_h_in_001_004+    86682.51997224252
Rh001_052_004-    i_052    tia_h_in_001_004-    121694.95973977765
Rh001_053_004+    i_053    tia_h_in_001_004+    120467.23948083716
Rh001_053_004-    i_053    tia_h_in_001_004-    82911.58654518423
Rh001_054_004+    i_054    tia_h_in_001_004+    71016.86155719089
Rh001_054_004-    i_054    tia_h_in_001_004-    118435.6276485873
Rh001_055_004+    i_055    tia_h_in_001_004+    120555.98373651963
Rh001_055_004-    i_055    tia_h_in_001_004-    81577.57650509985
Rh001_056_004+    i_056    tia_h_in_001_004+    118909.8920850459
Rh001_056_004-    i_056    tia_h_in_001_004-    59309.89476727268
Rh001_057_004+    i_057    tia_h_in_001_004+    121014.020332073
Rh001_057_004-    i_057    tia_h_in_001_004-    91445.46156508403
Rh001_058_004+    i_058    tia_h_in_001_004+    120139.1346020873
Rh001_058_004-    i_058    tia_h_in_001_004-    5000
Rh001_059_004+    i_059    tia_h_in_001_004+    120000
Rh001_059_004-    i_059    tia_h_in_001_004-    82730.24710319907
Rh001_060_004+    i_060    tia_h_in_001_004+    119015.64520998271
Rh001_060_004-    i_060    tia_h_in_001_004-    53374.69868048316
Rh001_061_004+    i_061    tia_h_in_001_004+    73039.51963163506
Rh001_061_004-    i_061    tia_h_in_001_004-    120858.42992084932
Rh001_062_004+    i_062    tia_h_in_001_004+    120000
Rh001_062_004-    i_062    tia_h_in_001_004-    60730.713376857566
Rh001_063_004+    i_063    tia_h_in_001_004+    77376.01064514743
Rh001_063_004-    i_063    tia_h_in_001_004-    121273.93777831194
Rh001_064_004+    i_064    tia_h_in_001_004+    81125.11964781997
Rh001_064_004-    i_064    tia_h_in_001_004-    120689.42380894619

* Neuron 5
Rh001_001_005+    i_001    tia_h_in_001_005+    119081.62861230587
Rh001_001_005-    i_001    tia_h_in_001_005-    23837.026895967017
Rh001_002_005+    i_002    tia_h_in_001_005+    119989.10230967081
Rh001_002_005-    i_002    tia_h_in_001_005-    120000
Rh001_003_005+    i_003    tia_h_in_001_005+    119882.3489619508
Rh001_003_005-    i_003    tia_h_in_001_005-    55971.00736380814
Rh001_004_005+    i_004    tia_h_in_001_005+    118388.72057933128
Rh001_004_005-    i_004    tia_h_in_001_005-    41988.25186154605
Rh001_005_005+    i_005    tia_h_in_001_005+    120035.89021907972
Rh001_005_005-    i_005    tia_h_in_001_005-    5000
Rh001_006_005+    i_006    tia_h_in_001_005+    111014.6853305869
Rh001_006_005-    i_006    tia_h_in_001_005-    121630.37064792066
Rh001_007_005+    i_007    tia_h_in_001_005+    121066.27698145871
Rh001_007_005-    i_007    tia_h_in_001_005-    45714.536379718826
Rh001_008_005+    i_008    tia_h_in_001_005+    120428.86874263959
Rh001_008_005-    i_008    tia_h_in_001_005-    82632.07598931543
Rh001_009_005+    i_009    tia_h_in_001_005+    92394.48061623196
Rh001_009_005-    i_009    tia_h_in_001_005-    118389.10413714605
Rh001_010_005+    i_010    tia_h_in_001_005+    23165.616657227656
Rh001_010_005-    i_010    tia_h_in_001_005-    120000
Rh001_011_005+    i_011    tia_h_in_001_005+    5000
Rh001_011_005-    i_011    tia_h_in_001_005-    121221.8698777941
Rh001_012_005+    i_012    tia_h_in_001_005+    90071.12313408803
Rh001_012_005-    i_012    tia_h_in_001_005-    120000
Rh001_013_005+    i_013    tia_h_in_001_005+    56804.731517626446
Rh001_013_005-    i_013    tia_h_in_001_005-    118947.52674911598
Rh001_014_005+    i_014    tia_h_in_001_005+    36042.88531694036
Rh001_014_005-    i_014    tia_h_in_001_005-    121284.58992499221
Rh001_015_005+    i_015    tia_h_in_001_005+    37687.19816426252
Rh001_015_005-    i_015    tia_h_in_001_005-    120000
Rh001_016_005+    i_016    tia_h_in_001_005+    42153.04563653967
Rh001_016_005-    i_016    tia_h_in_001_005-    120085.38242342469
Rh001_017_005+    i_017    tia_h_in_001_005+    120517.12263024448
Rh001_017_005-    i_017    tia_h_in_001_005-    85514.0027148246
Rh001_018_005+    i_018    tia_h_in_001_005+    120740.81897549669
Rh001_018_005-    i_018    tia_h_in_001_005-    72149.24572705936
Rh001_019_005+    i_019    tia_h_in_001_005+    42374.986432320315
Rh001_019_005-    i_019    tia_h_in_001_005-    119635.337975872
Rh001_020_005+    i_020    tia_h_in_001_005+    117181.25666244233
Rh001_020_005-    i_020    tia_h_in_001_005-    120000
Rh001_021_005+    i_021    tia_h_in_001_005+    121253.038338044
Rh001_021_005-    i_021    tia_h_in_001_005-    67783.92883589625
Rh001_022_005+    i_022    tia_h_in_001_005+    120823.86732302749
Rh001_022_005-    i_022    tia_h_in_001_005-    39175.459958698644
Rh001_023_005+    i_023    tia_h_in_001_005+    120590.2248021233
Rh001_023_005-    i_023    tia_h_in_001_005-    43734.614930267904
Rh001_024_005+    i_024    tia_h_in_001_005+    77555.72892692036
Rh001_024_005-    i_024    tia_h_in_001_005-    119218.73889756855
Rh001_025_005+    i_025    tia_h_in_001_005+    115957.52293858868
Rh001_025_005-    i_025    tia_h_in_001_005-    120473.57239866065
Rh001_026_005+    i_026    tia_h_in_001_005+    72555.83918695462
Rh001_026_005-    i_026    tia_h_in_001_005-    120131.21167054473
Rh001_027_005+    i_027    tia_h_in_001_005+    72622.81208641497
Rh001_027_005-    i_027    tia_h_in_001_005-    118809.95180087879
Rh001_028_005+    i_028    tia_h_in_001_005+    62586.47234876274
Rh001_028_005-    i_028    tia_h_in_001_005-    119049.07080184974
Rh001_029_005+    i_029    tia_h_in_001_005+    121693.06695810451
Rh001_029_005-    i_029    tia_h_in_001_005-    89622.05240674065
Rh001_030_005+    i_030    tia_h_in_001_005+    120805.88706966859
Rh001_030_005-    i_030    tia_h_in_001_005-    50242.2954857944
Rh001_031_005+    i_031    tia_h_in_001_005+    66935.4958721028
Rh001_031_005-    i_031    tia_h_in_001_005-    119649.94102496777
Rh001_032_005+    i_032    tia_h_in_001_005+    5000
Rh001_032_005-    i_032    tia_h_in_001_005-    120000
Rh001_033_005+    i_033    tia_h_in_001_005+    119216.07317519862
Rh001_033_005-    i_033    tia_h_in_001_005-    63880.13519789228
Rh001_034_005+    i_034    tia_h_in_001_005+    119884.70259494732
Rh001_034_005-    i_034    tia_h_in_001_005-    5000
Rh001_035_005+    i_035    tia_h_in_001_005+    119753.21043649327
Rh001_035_005-    i_035    tia_h_in_001_005-    71130.57851274888
Rh001_036_005+    i_036    tia_h_in_001_005+    108443.04166981769
Rh001_036_005-    i_036    tia_h_in_001_005-    120524.31195548935
Rh001_037_005+    i_037    tia_h_in_001_005+    113382.57857036505
Rh001_037_005-    i_037    tia_h_in_001_005-    119174.30997333945
Rh001_038_005+    i_038    tia_h_in_001_005+    118593.12640386481
Rh001_038_005-    i_038    tia_h_in_001_005-    78359.19362990253
Rh001_039_005+    i_039    tia_h_in_001_005+    120829.52117891195
Rh001_039_005-    i_039    tia_h_in_001_005-    60534.0038823434
Rh001_040_005+    i_040    tia_h_in_001_005+    79436.99809051339
Rh001_040_005-    i_040    tia_h_in_001_005-    5000
Rh001_041_005+    i_041    tia_h_in_001_005+    5000
Rh001_041_005-    i_041    tia_h_in_001_005-    120214.23127277866
Rh001_042_005+    i_042    tia_h_in_001_005+    119955.64173366713
Rh001_042_005-    i_042    tia_h_in_001_005-    81075.0743084
Rh001_043_005+    i_043    tia_h_in_001_005+    120477.54227571907
Rh001_043_005-    i_043    tia_h_in_001_005-    27791.750384357227
Rh001_044_005+    i_044    tia_h_in_001_005+    52868.45130629385
Rh001_044_005-    i_044    tia_h_in_001_005-    120945.02058511316
Rh001_045_005+    i_045    tia_h_in_001_005+    43407.43130374721
Rh001_045_005-    i_045    tia_h_in_001_005-    120600.42348727438
Rh001_046_005+    i_046    tia_h_in_001_005+    5000
Rh001_046_005-    i_046    tia_h_in_001_005-    89091.69693047366
Rh001_047_005+    i_047    tia_h_in_001_005+    118931.7706740132
Rh001_047_005-    i_047    tia_h_in_001_005-    28941.646157801133
Rh001_048_005+    i_048    tia_h_in_001_005+    119477.86904624088
Rh001_048_005-    i_048    tia_h_in_001_005-    49212.405936651536
Rh001_049_005+    i_049    tia_h_in_001_005+    120766.83721545826
Rh001_049_005-    i_049    tia_h_in_001_005-    96552.90544083864
Rh001_050_005+    i_050    tia_h_in_001_005+    96732.82398384079
Rh001_050_005-    i_050    tia_h_in_001_005-    120000
Rh001_051_005+    i_051    tia_h_in_001_005+    60053.49468682718
Rh001_051_005-    i_051    tia_h_in_001_005-    118628.68527463319
Rh001_052_005+    i_052    tia_h_in_001_005+    118897.95349659814
Rh001_052_005-    i_052    tia_h_in_001_005-    47912.01643821016
Rh001_053_005+    i_053    tia_h_in_001_005+    120000
Rh001_053_005-    i_053    tia_h_in_001_005-    122815.42284900161
Rh001_054_005+    i_054    tia_h_in_001_005+    41834.3732067741
Rh001_054_005-    i_054    tia_h_in_001_005-    121056.29543597491
Rh001_055_005+    i_055    tia_h_in_001_005+    38218.1755872526
Rh001_055_005-    i_055    tia_h_in_001_005-    121115.78866618275
Rh001_056_005+    i_056    tia_h_in_001_005+    120274.32981567425
Rh001_056_005-    i_056    tia_h_in_001_005-    54518.97693243147
Rh001_057_005+    i_057    tia_h_in_001_005+    58960.272812885916
Rh001_057_005-    i_057    tia_h_in_001_005-    120137.66096122412
Rh001_058_005+    i_058    tia_h_in_001_005+    120000
Rh001_058_005-    i_058    tia_h_in_001_005-    5000
Rh001_059_005+    i_059    tia_h_in_001_005+    64677.74516890222
Rh001_059_005-    i_059    tia_h_in_001_005-    120660.25386147355
Rh001_060_005+    i_060    tia_h_in_001_005+    103122.43342197071
Rh001_060_005-    i_060    tia_h_in_001_005-    121312.54789087342
Rh001_061_005+    i_061    tia_h_in_001_005+    119997.157069078
Rh001_061_005-    i_061    tia_h_in_001_005-    59873.11858722295
Rh001_062_005+    i_062    tia_h_in_001_005+    66728.99713229529
Rh001_062_005-    i_062    tia_h_in_001_005-    120985.46361924314
Rh001_063_005+    i_063    tia_h_in_001_005+    28283.637364233207
Rh001_063_005-    i_063    tia_h_in_001_005-    119067.25030230678
Rh001_064_005+    i_064    tia_h_in_001_005+    120150.26116462395
Rh001_064_005-    i_064    tia_h_in_001_005-    33769.095848337514

* Neuron 6
Rh001_001_006+    i_001    tia_h_in_001_006+    119936.8487415449
Rh001_001_006-    i_001    tia_h_in_001_006-    65502.860968724235
Rh001_002_006+    i_002    tia_h_in_001_006+    118912.16459258924
Rh001_002_006-    i_002    tia_h_in_001_006-    57577.145098998575
Rh001_003_006+    i_003    tia_h_in_001_006+    119762.81702186479
Rh001_003_006-    i_003    tia_h_in_001_006-    61954.52933900426
Rh001_004_006+    i_004    tia_h_in_001_006+    120275.6088722769
Rh001_004_006-    i_004    tia_h_in_001_006-    52389.057605756425
Rh001_005_006+    i_005    tia_h_in_001_006+    118968.38167560475
Rh001_005_006-    i_005    tia_h_in_001_006-    58709.520066739424
Rh001_006_006+    i_006    tia_h_in_001_006+    121699.50929533204
Rh001_006_006-    i_006    tia_h_in_001_006-    86164.50737406466
Rh001_007_006+    i_007    tia_h_in_001_006+    120000
Rh001_007_006-    i_007    tia_h_in_001_006-    120419.56785098833
Rh001_008_006+    i_008    tia_h_in_001_006+    5000
Rh001_008_006-    i_008    tia_h_in_001_006-    120180.16815326296
Rh001_009_006+    i_009    tia_h_in_001_006+    120275.73987664233
Rh001_009_006-    i_009    tia_h_in_001_006-    60415.508346633396
Rh001_010_006+    i_010    tia_h_in_001_006+    119930.80162399558
Rh001_010_006-    i_010    tia_h_in_001_006-    57880.08498225079
Rh001_011_006+    i_011    tia_h_in_001_006+    77467.37475101715
Rh001_011_006-    i_011    tia_h_in_001_006-    118979.30145477876
Rh001_012_006+    i_012    tia_h_in_001_006+    122027.70529307282
Rh001_012_006-    i_012    tia_h_in_001_006-    59723.92308190425
Rh001_013_006+    i_013    tia_h_in_001_006+    119810.01983823162
Rh001_013_006-    i_013    tia_h_in_001_006-    96783.75958372322
Rh001_014_006+    i_014    tia_h_in_001_006+    78477.59077038798
Rh001_014_006-    i_014    tia_h_in_001_006-    5000
Rh001_015_006+    i_015    tia_h_in_001_006+    120642.40424399747
Rh001_015_006-    i_015    tia_h_in_001_006-    73106.18070495175
Rh001_016_006+    i_016    tia_h_in_001_006+    119158.1283102575
Rh001_016_006-    i_016    tia_h_in_001_006-    101102.76405909797
Rh001_017_006+    i_017    tia_h_in_001_006+    119330.27081727436
Rh001_017_006-    i_017    tia_h_in_001_006-    103897.58320593425
Rh001_018_006+    i_018    tia_h_in_001_006+    120443.68268075302
Rh001_018_006-    i_018    tia_h_in_001_006-    87929.78131014785
Rh001_019_006+    i_019    tia_h_in_001_006+    122331.7974445496
Rh001_019_006-    i_019    tia_h_in_001_006-    70225.37991853981
Rh001_020_006+    i_020    tia_h_in_001_006+    118499.58659416744
Rh001_020_006-    i_020    tia_h_in_001_006-    54284.324209871644
Rh001_021_006+    i_021    tia_h_in_001_006+    118887.37925270315
Rh001_021_006-    i_021    tia_h_in_001_006-    57775.037888622785
Rh001_022_006+    i_022    tia_h_in_001_006+    120270.12903261934
Rh001_022_006-    i_022    tia_h_in_001_006-    69123.6662666779
Rh001_023_006+    i_023    tia_h_in_001_006+    55871.46634666341
Rh001_023_006-    i_023    tia_h_in_001_006-    120720.94593045492
Rh001_024_006+    i_024    tia_h_in_001_006+    121540.21705298289
Rh001_024_006-    i_024    tia_h_in_001_006-    72360.15623429476
Rh001_025_006+    i_025    tia_h_in_001_006+    121036.79147956193
Rh001_025_006-    i_025    tia_h_in_001_006-    63830.19291532338
Rh001_026_006+    i_026    tia_h_in_001_006+    95887.78232540577
Rh001_026_006-    i_026    tia_h_in_001_006-    120027.02222258307
Rh001_027_006+    i_027    tia_h_in_001_006+    94388.22564617706
Rh001_027_006-    i_027    tia_h_in_001_006-    119745.63765164258
Rh001_028_006+    i_028    tia_h_in_001_006+    74015.71756210613
Rh001_028_006-    i_028    tia_h_in_001_006-    119610.60659868324
Rh001_029_006+    i_029    tia_h_in_001_006+    63525.040704753774
Rh001_029_006-    i_029    tia_h_in_001_006-    119258.78354070603
Rh001_030_006+    i_030    tia_h_in_001_006+    72314.07465102863
Rh001_030_006-    i_030    tia_h_in_001_006-    119896.22721128086
Rh001_031_006+    i_031    tia_h_in_001_006+    119675.10166513316
Rh001_031_006-    i_031    tia_h_in_001_006-    51438.49380732103
Rh001_032_006+    i_032    tia_h_in_001_006+    113384.27492562086
Rh001_032_006-    i_032    tia_h_in_001_006-    119938.74707790189
Rh001_033_006+    i_033    tia_h_in_001_006+    69756.33998692186
Rh001_033_006-    i_033    tia_h_in_001_006-    120981.72074851883
Rh001_034_006+    i_034    tia_h_in_001_006+    120976.59584020243
Rh001_034_006-    i_034    tia_h_in_001_006-    99592.6159992284
Rh001_035_006+    i_035    tia_h_in_001_006+    120396.95090972052
Rh001_035_006-    i_035    tia_h_in_001_006-    66038.46900388246
Rh001_036_006+    i_036    tia_h_in_001_006+    55762.04012548326
Rh001_036_006-    i_036    tia_h_in_001_006-    120962.57891192076
Rh001_037_006+    i_037    tia_h_in_001_006+    120098.69886231392
Rh001_037_006-    i_037    tia_h_in_001_006-    75928.56164047107
Rh001_038_006+    i_038    tia_h_in_001_006+    118133.17644893665
Rh001_038_006-    i_038    tia_h_in_001_006-    67551.40689862249
Rh001_039_006+    i_039    tia_h_in_001_006+    120982.07261741812
Rh001_039_006-    i_039    tia_h_in_001_006-    55069.111595573704
Rh001_040_006+    i_040    tia_h_in_001_006+    120098.20497367381
Rh001_040_006-    i_040    tia_h_in_001_006-    120747.69978044633
Rh001_041_006+    i_041    tia_h_in_001_006+    81208.98245651954
Rh001_041_006-    i_041    tia_h_in_001_006-    121097.75454819702
Rh001_042_006+    i_042    tia_h_in_001_006+    99893.82443382672
Rh001_042_006-    i_042    tia_h_in_001_006-    119338.20095530919
Rh001_043_006+    i_043    tia_h_in_001_006+    120000
Rh001_043_006-    i_043    tia_h_in_001_006-    120355.40335500309
Rh001_044_006+    i_044    tia_h_in_001_006+    120722.1427872447
Rh001_044_006-    i_044    tia_h_in_001_006-    59635.377958927515
Rh001_045_006+    i_045    tia_h_in_001_006+    121168.35377099988
Rh001_045_006-    i_045    tia_h_in_001_006-    53741.60872893412
Rh001_046_006+    i_046    tia_h_in_001_006+    119638.81348315353
Rh001_046_006-    i_046    tia_h_in_001_006-    114453.40823561313
Rh001_047_006+    i_047    tia_h_in_001_006+    57556.19517014096
Rh001_047_006-    i_047    tia_h_in_001_006-    5000
Rh001_048_006+    i_048    tia_h_in_001_006+    120000
Rh001_048_006-    i_048    tia_h_in_001_006-    119686.43135515648
Rh001_049_006+    i_049    tia_h_in_001_006+    122003.39946458835
Rh001_049_006-    i_049    tia_h_in_001_006-    66880.90034350767
Rh001_050_006+    i_050    tia_h_in_001_006+    118193.86205782386
Rh001_050_006-    i_050    tia_h_in_001_006-    99456.77055110427
Rh001_051_006+    i_051    tia_h_in_001_006+    120269.85969929433
Rh001_051_006-    i_051    tia_h_in_001_006-    60923.69688183276
Rh001_052_006+    i_052    tia_h_in_001_006+    120104.2498818678
Rh001_052_006-    i_052    tia_h_in_001_006-    71848.03266238754
Rh001_053_006+    i_053    tia_h_in_001_006+    105124.165977452
Rh001_053_006-    i_053    tia_h_in_001_006-    119895.9507505888
Rh001_054_006+    i_054    tia_h_in_001_006+    75411.47123256022
Rh001_054_006-    i_054    tia_h_in_001_006-    119471.6523700792
Rh001_055_006+    i_055    tia_h_in_001_006+    60201.999391565274
Rh001_055_006-    i_055    tia_h_in_001_006-    118899.22748076779
Rh001_056_006+    i_056    tia_h_in_001_006+    120046.40512554366
Rh001_056_006-    i_056    tia_h_in_001_006-    54619.89644148975
Rh001_057_006+    i_057    tia_h_in_001_006+    67492.4360749775
Rh001_057_006-    i_057    tia_h_in_001_006-    120795.53330964106
Rh001_058_006+    i_058    tia_h_in_001_006+    120119.23864276231
Rh001_058_006-    i_058    tia_h_in_001_006-    5000
Rh001_059_006+    i_059    tia_h_in_001_006+    120000
Rh001_059_006-    i_059    tia_h_in_001_006-    119791.96087452113
Rh001_060_006+    i_060    tia_h_in_001_006+    60590.075159637956
Rh001_060_006-    i_060    tia_h_in_001_006-    118622.42572302936
Rh001_061_006+    i_061    tia_h_in_001_006+    119788.86825030211
Rh001_061_006-    i_061    tia_h_in_001_006-    114456.48409066317
Rh001_062_006+    i_062    tia_h_in_001_006+    58787.02218923607
Rh001_062_006-    i_062    tia_h_in_001_006-    121964.88681810988
Rh001_063_006+    i_063    tia_h_in_001_006+    120975.81327284343
Rh001_063_006-    i_063    tia_h_in_001_006-    56057.82452586123
Rh001_064_006+    i_064    tia_h_in_001_006+    119065.90264199901
Rh001_064_006-    i_064    tia_h_in_001_006-    120000

* Neuron 7
Rh001_001_007+    i_001    tia_h_in_001_007+    59072.53380206985
Rh001_001_007-    i_001    tia_h_in_001_007-    120642.50147575415
Rh001_002_007+    i_002    tia_h_in_001_007+    5000
Rh001_002_007-    i_002    tia_h_in_001_007-    94067.30020422998
Rh001_003_007+    i_003    tia_h_in_001_007+    118396.15927068506
Rh001_003_007-    i_003    tia_h_in_001_007-    77496.8217542851
Rh001_004_007+    i_004    tia_h_in_001_007+    44672.903614426315
Rh001_004_007-    i_004    tia_h_in_001_007-    119084.7352353184
Rh001_005_007+    i_005    tia_h_in_001_007+    71719.65753306926
Rh001_005_007-    i_005    tia_h_in_001_007-    120299.79236093278
Rh001_006_007+    i_006    tia_h_in_001_007+    83513.44904241452
Rh001_006_007-    i_006    tia_h_in_001_007-    120142.85778961114
Rh001_007_007+    i_007    tia_h_in_001_007+    56850.872798444165
Rh001_007_007-    i_007    tia_h_in_001_007-    119931.6084283373
Rh001_008_007+    i_008    tia_h_in_001_007+    61525.09396513786
Rh001_008_007-    i_008    tia_h_in_001_007-    120205.2780213198
Rh001_009_007+    i_009    tia_h_in_001_007+    119937.20056394949
Rh001_009_007-    i_009    tia_h_in_001_007-    29093.46558298536
Rh001_010_007+    i_010    tia_h_in_001_007+    119917.04333061294
Rh001_010_007-    i_010    tia_h_in_001_007-    50211.58397446003
Rh001_011_007+    i_011    tia_h_in_001_007+    43711.10822936231
Rh001_011_007-    i_011    tia_h_in_001_007-    121474.20881588315
Rh001_012_007+    i_012    tia_h_in_001_007+    120000
Rh001_012_007-    i_012    tia_h_in_001_007-    119716.90118753022
Rh001_013_007+    i_013    tia_h_in_001_007+    118292.3109552282
Rh001_013_007-    i_013    tia_h_in_001_007-    120606.89632603475
Rh001_014_007+    i_014    tia_h_in_001_007+    42192.41954886613
Rh001_014_007-    i_014    tia_h_in_001_007-    120798.00282462058
Rh001_015_007+    i_015    tia_h_in_001_007+    80080.50783230223
Rh001_015_007-    i_015    tia_h_in_001_007-    120000
Rh001_016_007+    i_016    tia_h_in_001_007+    42065.82587112425
Rh001_016_007-    i_016    tia_h_in_001_007-    119540.26242752881
Rh001_017_007+    i_017    tia_h_in_001_007+    120021.75603665218
Rh001_017_007-    i_017    tia_h_in_001_007-    47881.1368331632
Rh001_018_007+    i_018    tia_h_in_001_007+    120000
Rh001_018_007-    i_018    tia_h_in_001_007-    53119.57470969745
Rh001_019_007+    i_019    tia_h_in_001_007+    5000
Rh001_019_007-    i_019    tia_h_in_001_007-    34658.318987538645
Rh001_020_007+    i_020    tia_h_in_001_007+    120511.04128388873
Rh001_020_007-    i_020    tia_h_in_001_007-    87552.76390431207
Rh001_021_007+    i_021    tia_h_in_001_007+    117306.83686615167
Rh001_021_007-    i_021    tia_h_in_001_007-    67293.6026922004
Rh001_022_007+    i_022    tia_h_in_001_007+    119615.2017995276
Rh001_022_007-    i_022    tia_h_in_001_007-    41371.290889594195
Rh001_023_007+    i_023    tia_h_in_001_007+    119243.49758837876
Rh001_023_007-    i_023    tia_h_in_001_007-    120000
Rh001_024_007+    i_024    tia_h_in_001_007+    101225.2917039336
Rh001_024_007-    i_024    tia_h_in_001_007-    120442.8947005236
Rh001_025_007+    i_025    tia_h_in_001_007+    65453.94677742859
Rh001_025_007-    i_025    tia_h_in_001_007-    5000
Rh001_026_007+    i_026    tia_h_in_001_007+    37591.16117389839
Rh001_026_007-    i_026    tia_h_in_001_007-    119674.45224039578
Rh001_027_007+    i_027    tia_h_in_001_007+    98181.21552270639
Rh001_027_007-    i_027    tia_h_in_001_007-    120177.21073985107
Rh001_028_007+    i_028    tia_h_in_001_007+    118730.44652629727
Rh001_028_007-    i_028    tia_h_in_001_007-    64914.58343226704
Rh001_029_007+    i_029    tia_h_in_001_007+    119367.85410553594
Rh001_029_007-    i_029    tia_h_in_001_007-    51811.5679697719
Rh001_030_007+    i_030    tia_h_in_001_007+    118193.86187128935
Rh001_030_007-    i_030    tia_h_in_001_007-    102446.59380548786
Rh001_031_007+    i_031    tia_h_in_001_007+    119673.62404881298
Rh001_031_007-    i_031    tia_h_in_001_007-    67226.86868629142
Rh001_032_007+    i_032    tia_h_in_001_007+    120747.90666448562
Rh001_032_007-    i_032    tia_h_in_001_007-    80177.40562856627
Rh001_033_007+    i_033    tia_h_in_001_007+    95077.14103370807
Rh001_033_007-    i_033    tia_h_in_001_007-    121397.3096552531
Rh001_034_007+    i_034    tia_h_in_001_007+    49380.493950856646
Rh001_034_007-    i_034    tia_h_in_001_007-    120479.02267686595
Rh001_035_007+    i_035    tia_h_in_001_007+    120000
Rh001_035_007-    i_035    tia_h_in_001_007-    31687.09929119376
Rh001_036_007+    i_036    tia_h_in_001_007+    5000
Rh001_036_007-    i_036    tia_h_in_001_007-    98647.94268364881
Rh001_037_007+    i_037    tia_h_in_001_007+    64361.92565175169
Rh001_037_007-    i_037    tia_h_in_001_007-    119698.22735958495
Rh001_038_007+    i_038    tia_h_in_001_007+    119144.16674485832
Rh001_038_007-    i_038    tia_h_in_001_007-    47722.343487772785
Rh001_039_007+    i_039    tia_h_in_001_007+    62012.689872985204
Rh001_039_007-    i_039    tia_h_in_001_007-    121700.35372593996
Rh001_040_007+    i_040    tia_h_in_001_007+    120373.74798266096
Rh001_040_007-    i_040    tia_h_in_001_007-    53482.918773990095
Rh001_041_007+    i_041    tia_h_in_001_007+    5000
Rh001_041_007-    i_041    tia_h_in_001_007-    121423.1033263421
Rh001_042_007+    i_042    tia_h_in_001_007+    57499.1062205748
Rh001_042_007-    i_042    tia_h_in_001_007-    121564.63348998757
Rh001_043_007+    i_043    tia_h_in_001_007+    120974.34280371829
Rh001_043_007-    i_043    tia_h_in_001_007-    5000
Rh001_044_007+    i_044    tia_h_in_001_007+    87582.7840485022
Rh001_044_007-    i_044    tia_h_in_001_007-    120164.53854027795
Rh001_045_007+    i_045    tia_h_in_001_007+    120805.08301430685
Rh001_045_007-    i_045    tia_h_in_001_007-    39158.81177857194
Rh001_046_007+    i_046    tia_h_in_001_007+    108971.06747178978
Rh001_046_007-    i_046    tia_h_in_001_007-    5000
Rh001_047_007+    i_047    tia_h_in_001_007+    49231.83012613928
Rh001_047_007-    i_047    tia_h_in_001_007-    5000
Rh001_048_007+    i_048    tia_h_in_001_007+    79560.16460716736
Rh001_048_007-    i_048    tia_h_in_001_007-    120232.55382223867
Rh001_049_007+    i_049    tia_h_in_001_007+    5000
Rh001_049_007-    i_049    tia_h_in_001_007-    118777.6353110569
Rh001_050_007+    i_050    tia_h_in_001_007+    82050.70090991548
Rh001_050_007-    i_050    tia_h_in_001_007-    119667.7138709335
Rh001_051_007+    i_051    tia_h_in_001_007+    30768.317887666446
Rh001_051_007-    i_051    tia_h_in_001_007-    119423.49699705327
Rh001_052_007+    i_052    tia_h_in_001_007+    120000
Rh001_052_007-    i_052    tia_h_in_001_007-    119142.98194016104
Rh001_053_007+    i_053    tia_h_in_001_007+    38446.3131124895
Rh001_053_007-    i_053    tia_h_in_001_007-    119749.003463634
Rh001_054_007+    i_054    tia_h_in_001_007+    23930.224210493405
Rh001_054_007-    i_054    tia_h_in_001_007-    120622.39706198713
Rh001_055_007+    i_055    tia_h_in_001_007+    34905.292058333755
Rh001_055_007-    i_055    tia_h_in_001_007-    121104.34090124191
Rh001_056_007+    i_056    tia_h_in_001_007+    53965.86125950682
Rh001_056_007-    i_056    tia_h_in_001_007-    121702.0035930592
Rh001_057_007+    i_057    tia_h_in_001_007+    61384.18384710241
Rh001_057_007-    i_057    tia_h_in_001_007-    120000
Rh001_058_007+    i_058    tia_h_in_001_007+    121019.16847555892
Rh001_058_007-    i_058    tia_h_in_001_007-    72073.34252442692
Rh001_059_007+    i_059    tia_h_in_001_007+    119330.01608273109
Rh001_059_007-    i_059    tia_h_in_001_007-    43175.438880788155
Rh001_060_007+    i_060    tia_h_in_001_007+    119487.17156285931
Rh001_060_007-    i_060    tia_h_in_001_007-    120000
Rh001_061_007+    i_061    tia_h_in_001_007+    63651.600125597426
Rh001_061_007-    i_061    tia_h_in_001_007-    119306.28111545042
Rh001_062_007+    i_062    tia_h_in_001_007+    120000
Rh001_062_007-    i_062    tia_h_in_001_007-    22428.326783631284
Rh001_063_007+    i_063    tia_h_in_001_007+    120000
Rh001_063_007-    i_063    tia_h_in_001_007-    17812.3686341136
Rh001_064_007+    i_064    tia_h_in_001_007+    118552.20384167683
Rh001_064_007-    i_064    tia_h_in_001_007-    5000

* Neuron 8
Rh001_001_008+    i_001    tia_h_in_001_008+    118866.14374425636
Rh001_001_008-    i_001    tia_h_in_001_008-    39600.900576564774
Rh001_002_008+    i_002    tia_h_in_001_008+    45365.35973811732
Rh001_002_008-    i_002    tia_h_in_001_008-    117804.16013707081
Rh001_003_008+    i_003    tia_h_in_001_008+    119596.89149027616
Rh001_003_008-    i_003    tia_h_in_001_008-    56502.454495203674
Rh001_004_008+    i_004    tia_h_in_001_008+    120000
Rh001_004_008-    i_004    tia_h_in_001_008-    71456.57657061938
Rh001_005_008+    i_005    tia_h_in_001_008+    107406.63888247861
Rh001_005_008-    i_005    tia_h_in_001_008-    120022.33786089848
Rh001_006_008+    i_006    tia_h_in_001_008+    51554.84649376765
Rh001_006_008-    i_006    tia_h_in_001_008-    119961.69906228142
Rh001_007_008+    i_007    tia_h_in_001_008+    83155.40328962315
Rh001_007_008-    i_007    tia_h_in_001_008-    120948.44445417791
Rh001_008_008+    i_008    tia_h_in_001_008+    31784.304620175757
Rh001_008_008-    i_008    tia_h_in_001_008-    120439.65896761017
Rh001_009_008+    i_009    tia_h_in_001_008+    71168.65055190744
Rh001_009_008-    i_009    tia_h_in_001_008-    118324.00713151903
Rh001_010_008+    i_010    tia_h_in_001_008+    85751.56312323849
Rh001_010_008-    i_010    tia_h_in_001_008-    120667.49355623001
Rh001_011_008+    i_011    tia_h_in_001_008+    48649.83845051985
Rh001_011_008-    i_011    tia_h_in_001_008-    120859.83964857884
Rh001_012_008+    i_012    tia_h_in_001_008+    119746.90407087478
Rh001_012_008-    i_012    tia_h_in_001_008-    31987.239626890805
Rh001_013_008+    i_013    tia_h_in_001_008+    119595.18349329123
Rh001_013_008-    i_013    tia_h_in_001_008-    81923.71429546317
Rh001_014_008+    i_014    tia_h_in_001_008+    118999.89327620181
Rh001_014_008-    i_014    tia_h_in_001_008-    49281.56504044414
Rh001_015_008+    i_015    tia_h_in_001_008+    120093.73465868672
Rh001_015_008-    i_015    tia_h_in_001_008-    120000
Rh001_016_008+    i_016    tia_h_in_001_008+    121245.78369243586
Rh001_016_008-    i_016    tia_h_in_001_008-    95324.83144651742
Rh001_017_008+    i_017    tia_h_in_001_008+    32380.413680867023
Rh001_017_008-    i_017    tia_h_in_001_008-    119012.4119979256
Rh001_018_008+    i_018    tia_h_in_001_008+    56023.7892947411
Rh001_018_008-    i_018    tia_h_in_001_008-    119758.19472551913
Rh001_019_008+    i_019    tia_h_in_001_008+    33232.6488144573
Rh001_019_008-    i_019    tia_h_in_001_008-    119777.68681742686
Rh001_020_008+    i_020    tia_h_in_001_008+    31484.619456086115
Rh001_020_008-    i_020    tia_h_in_001_008-    119631.26879024718
Rh001_021_008+    i_021    tia_h_in_001_008+    60401.64861949993
Rh001_021_008-    i_021    tia_h_in_001_008-    121037.03145431267
Rh001_022_008+    i_022    tia_h_in_001_008+    121630.7910631755
Rh001_022_008-    i_022    tia_h_in_001_008-    48606.587257821986
Rh001_023_008+    i_023    tia_h_in_001_008+    92732.92249967669
Rh001_023_008-    i_023    tia_h_in_001_008-    120000
Rh001_024_008+    i_024    tia_h_in_001_008+    119577.7504295201
Rh001_024_008-    i_024    tia_h_in_001_008-    29195.389295556957
Rh001_025_008+    i_025    tia_h_in_001_008+    111019.64042759
Rh001_025_008-    i_025    tia_h_in_001_008-    119333.17262488585
Rh001_026_008+    i_026    tia_h_in_001_008+    120432.14826718812
Rh001_026_008-    i_026    tia_h_in_001_008-    57535.209585879325
Rh001_027_008+    i_027    tia_h_in_001_008+    79869.96974887834
Rh001_027_008-    i_027    tia_h_in_001_008-    119999.16681290038
Rh001_028_008+    i_028    tia_h_in_001_008+    39472.652102956046
Rh001_028_008-    i_028    tia_h_in_001_008-    120576.16182405861
Rh001_029_008+    i_029    tia_h_in_001_008+    121250.03352210642
Rh001_029_008-    i_029    tia_h_in_001_008-    88072.95353309077
Rh001_030_008+    i_030    tia_h_in_001_008+    119384.71198320485
Rh001_030_008-    i_030    tia_h_in_001_008-    113530.36306451829
Rh001_031_008+    i_031    tia_h_in_001_008+    118790.1996562059
Rh001_031_008-    i_031    tia_h_in_001_008-    120000
Rh001_032_008+    i_032    tia_h_in_001_008+    118786.73658638935
Rh001_032_008-    i_032    tia_h_in_001_008-    84356.22054040234
Rh001_033_008+    i_033    tia_h_in_001_008+    120636.34632825814
Rh001_033_008-    i_033    tia_h_in_001_008-    62316.19272873343
Rh001_034_008+    i_034    tia_h_in_001_008+    68002.87894594007
Rh001_034_008-    i_034    tia_h_in_001_008-    120000
Rh001_035_008+    i_035    tia_h_in_001_008+    91480.95714008682
Rh001_035_008-    i_035    tia_h_in_001_008-    121108.29224479514
Rh001_036_008+    i_036    tia_h_in_001_008+    119149.58033371824
Rh001_036_008-    i_036    tia_h_in_001_008-    35564.61890720878
Rh001_037_008+    i_037    tia_h_in_001_008+    55044.396343409215
Rh001_037_008-    i_037    tia_h_in_001_008-    120931.79092305816
Rh001_038_008+    i_038    tia_h_in_001_008+    50722.25952820306
Rh001_038_008-    i_038    tia_h_in_001_008-    120753.93444987164
Rh001_039_008+    i_039    tia_h_in_001_008+    118951.8324549659
Rh001_039_008-    i_039    tia_h_in_001_008-    110341.44185990778
Rh001_040_008+    i_040    tia_h_in_001_008+    47010.39208026604
Rh001_040_008-    i_040    tia_h_in_001_008-    120016.75150893503
Rh001_041_008+    i_041    tia_h_in_001_008+    121280.57337950772
Rh001_041_008-    i_041    tia_h_in_001_008-    56602.97490586507
Rh001_042_008+    i_042    tia_h_in_001_008+    120535.38633983566
Rh001_042_008-    i_042    tia_h_in_001_008-    32620.5455590458
Rh001_043_008+    i_043    tia_h_in_001_008+    119929.41193472967
Rh001_043_008-    i_043    tia_h_in_001_008-    49015.4338285898
Rh001_044_008+    i_044    tia_h_in_001_008+    121888.14548875522
Rh001_044_008-    i_044    tia_h_in_001_008-    45586.27185317038
Rh001_045_008+    i_045    tia_h_in_001_008+    82829.36900406948
Rh001_045_008-    i_045    tia_h_in_001_008-    121342.57507310995
Rh001_046_008+    i_046    tia_h_in_001_008+    34787.75811853994
Rh001_046_008-    i_046    tia_h_in_001_008-    119125.4012407887
Rh001_047_008+    i_047    tia_h_in_001_008+    55907.11299877083
Rh001_047_008-    i_047    tia_h_in_001_008-    120566.74537754344
Rh001_048_008+    i_048    tia_h_in_001_008+    24300.373544422608
Rh001_048_008-    i_048    tia_h_in_001_008-    118998.01445405492
Rh001_049_008+    i_049    tia_h_in_001_008+    120048.9217958316
Rh001_049_008-    i_049    tia_h_in_001_008-    68398.962890391
Rh001_050_008+    i_050    tia_h_in_001_008+    75340.82407405376
Rh001_050_008-    i_050    tia_h_in_001_008-    119458.47639009656
Rh001_051_008+    i_051    tia_h_in_001_008+    99435.69300808494
Rh001_051_008-    i_051    tia_h_in_001_008-    121717.17159251611
Rh001_052_008+    i_052    tia_h_in_001_008+    47665.518066181845
Rh001_052_008-    i_052    tia_h_in_001_008-    119247.35623903493
Rh001_053_008+    i_053    tia_h_in_001_008+    5000
Rh001_053_008-    i_053    tia_h_in_001_008-    118941.23260571202
Rh001_054_008+    i_054    tia_h_in_001_008+    31942.301896500303
Rh001_054_008-    i_054    tia_h_in_001_008-    120155.9780172134
Rh001_055_008+    i_055    tia_h_in_001_008+    27379.836303918382
Rh001_055_008-    i_055    tia_h_in_001_008-    122256.08779842338
Rh001_056_008+    i_056    tia_h_in_001_008+    67354.24510720062
Rh001_056_008-    i_056    tia_h_in_001_008-    118447.84358348792
Rh001_057_008+    i_057    tia_h_in_001_008+    121465.05308567252
Rh001_057_008-    i_057    tia_h_in_001_008-    99830.0522903742
Rh001_058_008+    i_058    tia_h_in_001_008+    119944.06454451605
Rh001_058_008-    i_058    tia_h_in_001_008-    77896.54995192509
Rh001_059_008+    i_059    tia_h_in_001_008+    88152.77859968797
Rh001_059_008-    i_059    tia_h_in_001_008-    119114.48598366922
Rh001_060_008+    i_060    tia_h_in_001_008+    119296.2261891149
Rh001_060_008-    i_060    tia_h_in_001_008-    22315.43556298645
Rh001_061_008+    i_061    tia_h_in_001_008+    120300.82280883982
Rh001_061_008-    i_061    tia_h_in_001_008-    36211.817432419106
Rh001_062_008+    i_062    tia_h_in_001_008+    120000
Rh001_062_008-    i_062    tia_h_in_001_008-    26101.202032580284
Rh001_063_008+    i_063    tia_h_in_001_008+    121225.36807084635
Rh001_063_008-    i_063    tia_h_in_001_008-    15550.120834907924
Rh001_064_008+    i_064    tia_h_in_001_008+    120802.48700791919
Rh001_064_008-    i_064    tia_h_in_001_008-    16213.669217334815

* Neuron 9
Rh001_001_009+    i_001    tia_h_in_001_009+    63706.9846044507
Rh001_001_009-    i_001    tia_h_in_001_009-    120000
Rh001_002_009+    i_002    tia_h_in_001_009+    118988.63656101757
Rh001_002_009-    i_002    tia_h_in_001_009-    38273.91175335973
Rh001_003_009+    i_003    tia_h_in_001_009+    120548.18405435706
Rh001_003_009-    i_003    tia_h_in_001_009-    82521.71440882212
Rh001_004_009+    i_004    tia_h_in_001_009+    80472.82399051049
Rh001_004_009-    i_004    tia_h_in_001_009-    120420.79456014212
Rh001_005_009+    i_005    tia_h_in_001_009+    103376.96107462981
Rh001_005_009-    i_005    tia_h_in_001_009-    119558.51837370823
Rh001_006_009+    i_006    tia_h_in_001_009+    64224.071823564664
Rh001_006_009-    i_006    tia_h_in_001_009-    119126.16072268625
Rh001_007_009+    i_007    tia_h_in_001_009+    120000
Rh001_007_009-    i_007    tia_h_in_001_009-    119971.73795186408
Rh001_008_009+    i_008    tia_h_in_001_009+    5000
Rh001_008_009-    i_008    tia_h_in_001_009-    120313.04765838341
Rh001_009_009+    i_009    tia_h_in_001_009+    5000
Rh001_009_009-    i_009    tia_h_in_001_009-    120200.63818609393
Rh001_010_009+    i_010    tia_h_in_001_009+    118777.51412002102
Rh001_010_009-    i_010    tia_h_in_001_009-    61197.62903415241
Rh001_011_009+    i_011    tia_h_in_001_009+    89669.89607352576
Rh001_011_009-    i_011    tia_h_in_001_009-    119226.11020793726
Rh001_012_009+    i_012    tia_h_in_001_009+    50412.86714480424
Rh001_012_009-    i_012    tia_h_in_001_009-    120570.31906716614
Rh001_013_009+    i_013    tia_h_in_001_009+    120285.7202231417
Rh001_013_009-    i_013    tia_h_in_001_009-    61209.77796448012
Rh001_014_009+    i_014    tia_h_in_001_009+    118769.179364206
Rh001_014_009-    i_014    tia_h_in_001_009-    120000
Rh001_015_009+    i_015    tia_h_in_001_009+    120878.86184874736
Rh001_015_009-    i_015    tia_h_in_001_009-    66509.85502150666
Rh001_016_009+    i_016    tia_h_in_001_009+    120218.79943046186
Rh001_016_009-    i_016    tia_h_in_001_009-    29790.665165982362
Rh001_017_009+    i_017    tia_h_in_001_009+    5000
Rh001_017_009-    i_017    tia_h_in_001_009-    120000
Rh001_018_009+    i_018    tia_h_in_001_009+    28592.776087236067
Rh001_018_009-    i_018    tia_h_in_001_009-    120310.37018474478
Rh001_019_009+    i_019    tia_h_in_001_009+    87835.46872373845
Rh001_019_009-    i_019    tia_h_in_001_009-    119834.606109384
Rh001_020_009+    i_020    tia_h_in_001_009+    119714.47422266136
Rh001_020_009-    i_020    tia_h_in_001_009-    86241.01839980221
Rh001_021_009+    i_021    tia_h_in_001_009+    120238.40131752203
Rh001_021_009-    i_021    tia_h_in_001_009-    50112.501339345734
Rh001_022_009+    i_022    tia_h_in_001_009+    120167.87717730328
Rh001_022_009-    i_022    tia_h_in_001_009-    5000
Rh001_023_009+    i_023    tia_h_in_001_009+    119943.47577961604
Rh001_023_009-    i_023    tia_h_in_001_009-    117714.88183209795
Rh001_024_009+    i_024    tia_h_in_001_009+    54095.88413696677
Rh001_024_009-    i_024    tia_h_in_001_009-    119526.05211998215
Rh001_025_009+    i_025    tia_h_in_001_009+    120269.10771081244
Rh001_025_009-    i_025    tia_h_in_001_009-    26287.740866058422
Rh001_026_009+    i_026    tia_h_in_001_009+    99947.44201164602
Rh001_026_009-    i_026    tia_h_in_001_009-    118423.10966898351
Rh001_027_009+    i_027    tia_h_in_001_009+    119635.17616244826
Rh001_027_009-    i_027    tia_h_in_001_009-    88104.07955968869
Rh001_028_009+    i_028    tia_h_in_001_009+    83864.54556146065
Rh001_028_009-    i_028    tia_h_in_001_009-    119167.36031166822
Rh001_029_009+    i_029    tia_h_in_001_009+    76970.3453017631
Rh001_029_009-    i_029    tia_h_in_001_009-    119302.00285239595
Rh001_030_009+    i_030    tia_h_in_001_009+    74601.73437818696
Rh001_030_009-    i_030    tia_h_in_001_009-    120682.67225460685
Rh001_031_009+    i_031    tia_h_in_001_009+    54198.3014377626
Rh001_031_009-    i_031    tia_h_in_001_009-    119217.43510791312
Rh001_032_009+    i_032    tia_h_in_001_009+    40932.995315042026
Rh001_032_009-    i_032    tia_h_in_001_009-    119950.3321479578
Rh001_033_009+    i_033    tia_h_in_001_009+    38465.763789839446
Rh001_033_009-    i_033    tia_h_in_001_009-    119783.49477852906
Rh001_034_009+    i_034    tia_h_in_001_009+    64342.73943489871
Rh001_034_009-    i_034    tia_h_in_001_009-    119791.48027667007
Rh001_035_009+    i_035    tia_h_in_001_009+    119547.40158993004
Rh001_035_009-    i_035    tia_h_in_001_009-    63165.80086452789
Rh001_036_009+    i_036    tia_h_in_001_009+    100463.82262801252
Rh001_036_009-    i_036    tia_h_in_001_009-    119952.71202480338
Rh001_037_009+    i_037    tia_h_in_001_009+    118373.24707555478
Rh001_037_009-    i_037    tia_h_in_001_009-    104492.52808504635
Rh001_038_009+    i_038    tia_h_in_001_009+    120000
Rh001_038_009-    i_038    tia_h_in_001_009-    119781.21005758853
Rh001_039_009+    i_039    tia_h_in_001_009+    120793.94485215441
Rh001_039_009-    i_039    tia_h_in_001_009-    5000
Rh001_040_009+    i_040    tia_h_in_001_009+    50388.5575367172
Rh001_040_009-    i_040    tia_h_in_001_009-    119511.64464785837
Rh001_041_009+    i_041    tia_h_in_001_009+    33577.23720955747
Rh001_041_009-    i_041    tia_h_in_001_009-    119462.93022804345
Rh001_042_009+    i_042    tia_h_in_001_009+    81433.4663729821
Rh001_042_009-    i_042    tia_h_in_001_009-    118950.32523946304
Rh001_043_009+    i_043    tia_h_in_001_009+    80806.75564632003
Rh001_043_009-    i_043    tia_h_in_001_009-    120716.88916918305
Rh001_044_009+    i_044    tia_h_in_001_009+    37361.49300571458
Rh001_044_009-    i_044    tia_h_in_001_009-    119293.9288929917
Rh001_045_009+    i_045    tia_h_in_001_009+    33248.59829972157
Rh001_045_009-    i_045    tia_h_in_001_009-    121747.60806518591
Rh001_046_009+    i_046    tia_h_in_001_009+    77278.48571701928
Rh001_046_009-    i_046    tia_h_in_001_009-    119298.08635861143
Rh001_047_009+    i_047    tia_h_in_001_009+    40919.34447591468
Rh001_047_009-    i_047    tia_h_in_001_009-    5000
Rh001_048_009+    i_048    tia_h_in_001_009+    24173.065637132266
Rh001_048_009-    i_048    tia_h_in_001_009-    119634.4559032895
Rh001_049_009+    i_049    tia_h_in_001_009+    120735.01967267162
Rh001_049_009-    i_049    tia_h_in_001_009-    86145.69971511261
Rh001_050_009+    i_050    tia_h_in_001_009+    78545.73528359615
Rh001_050_009-    i_050    tia_h_in_001_009-    120688.32870958744
Rh001_051_009+    i_051    tia_h_in_001_009+    120295.74351733582
Rh001_051_009-    i_051    tia_h_in_001_009-    37306.70692836042
Rh001_052_009+    i_052    tia_h_in_001_009+    120000
Rh001_052_009-    i_052    tia_h_in_001_009-    84779.10242493609
Rh001_053_009+    i_053    tia_h_in_001_009+    5000
Rh001_053_009-    i_053    tia_h_in_001_009-    52123.16279331561
Rh001_054_009+    i_054    tia_h_in_001_009+    121063.48419519835
Rh001_054_009-    i_054    tia_h_in_001_009-    114547.1780033869
Rh001_055_009+    i_055    tia_h_in_001_009+    49961.283451071606
Rh001_055_009-    i_055    tia_h_in_001_009-    119954.79592986211
Rh001_056_009+    i_056    tia_h_in_001_009+    119290.67056028335
Rh001_056_009-    i_056    tia_h_in_001_009-    45432.34339225255
Rh001_057_009+    i_057    tia_h_in_001_009+    119538.03017894085
Rh001_057_009-    i_057    tia_h_in_001_009-    54474.9146720373
Rh001_058_009+    i_058    tia_h_in_001_009+    119228.48324750035
Rh001_058_009-    i_058    tia_h_in_001_009-    48185.23025297832
Rh001_059_009+    i_059    tia_h_in_001_009+    76965.3980167635
Rh001_059_009-    i_059    tia_h_in_001_009-    119445.99577422206
Rh001_060_009+    i_060    tia_h_in_001_009+    119857.44357729777
Rh001_060_009-    i_060    tia_h_in_001_009-    47603.24165043898
Rh001_061_009+    i_061    tia_h_in_001_009+    121785.22960181124
Rh001_061_009-    i_061    tia_h_in_001_009-    35771.98891459064
Rh001_062_009+    i_062    tia_h_in_001_009+    119643.51719524025
Rh001_062_009-    i_062    tia_h_in_001_009-    53331.901515770995
Rh001_063_009+    i_063    tia_h_in_001_009+    120389.67356485328
Rh001_063_009-    i_063    tia_h_in_001_009-    21156.038309369498
Rh001_064_009+    i_064    tia_h_in_001_009+    119371.60997037319
Rh001_064_009-    i_064    tia_h_in_001_009-    14672.443760823315

* Neuron 10
Rh001_001_010+    i_001    tia_h_in_001_010+    69669.83863805435
Rh001_001_010-    i_001    tia_h_in_001_010-    119677.2557145131
Rh001_002_010+    i_002    tia_h_in_001_010+    119701.60252639808
Rh001_002_010-    i_002    tia_h_in_001_010-    56597.51457478093
Rh001_003_010+    i_003    tia_h_in_001_010+    108181.39386861172
Rh001_003_010-    i_003    tia_h_in_001_010-    121263.05791545204
Rh001_004_010+    i_004    tia_h_in_001_010+    58019.30803762199
Rh001_004_010-    i_004    tia_h_in_001_010-    117982.29571741969
Rh001_005_010+    i_005    tia_h_in_001_010+    101868.47362900521
Rh001_005_010-    i_005    tia_h_in_001_010-    118711.34796576081
Rh001_006_010+    i_006    tia_h_in_001_010+    93063.87122435485
Rh001_006_010-    i_006    tia_h_in_001_010-    120638.08560297257
Rh001_007_010+    i_007    tia_h_in_001_010+    118659.18665808305
Rh001_007_010-    i_007    tia_h_in_001_010-    67730.47765333671
Rh001_008_010+    i_008    tia_h_in_001_010+    119806.76737735921
Rh001_008_010-    i_008    tia_h_in_001_010-    113363.12762467621
Rh001_009_010+    i_009    tia_h_in_001_010+    119537.89571959297
Rh001_009_010-    i_009    tia_h_in_001_010-    119637.55570348528
Rh001_010_010+    i_010    tia_h_in_001_010+    94420.34065486227
Rh001_010_010-    i_010    tia_h_in_001_010-    120440.16415181877
Rh001_011_010+    i_011    tia_h_in_001_010+    5000
Rh001_011_010-    i_011    tia_h_in_001_010-    121198.36222134758
Rh001_012_010+    i_012    tia_h_in_001_010+    59117.908196857876
Rh001_012_010-    i_012    tia_h_in_001_010-    119417.1838275226
Rh001_013_010+    i_013    tia_h_in_001_010+    120290.0307758832
Rh001_013_010-    i_013    tia_h_in_001_010-    60533.258899259126
Rh001_014_010+    i_014    tia_h_in_001_010+    5000
Rh001_014_010-    i_014    tia_h_in_001_010-    119425.45824262092
Rh001_015_010+    i_015    tia_h_in_001_010+    118178.23586354606
Rh001_015_010-    i_015    tia_h_in_001_010-    120000
Rh001_016_010+    i_016    tia_h_in_001_010+    120746.77771673493
Rh001_016_010-    i_016    tia_h_in_001_010-    59480.840126303105
Rh001_017_010+    i_017    tia_h_in_001_010+    120839.84757746209
Rh001_017_010-    i_017    tia_h_in_001_010-    103944.62929316428
Rh001_018_010+    i_018    tia_h_in_001_010+    119998.63395714336
Rh001_018_010-    i_018    tia_h_in_001_010-    55863.05995493351
Rh001_019_010+    i_019    tia_h_in_001_010+    67125.67229642904
Rh001_019_010-    i_019    tia_h_in_001_010-    120298.82349980398
Rh001_020_010+    i_020    tia_h_in_001_010+    109672.13599703941
Rh001_020_010-    i_020    tia_h_in_001_010-    119799.99591489612
Rh001_021_010+    i_021    tia_h_in_001_010+    118919.53487191584
Rh001_021_010-    i_021    tia_h_in_001_010-    69988.26254710525
Rh001_022_010+    i_022    tia_h_in_001_010+    73889.74779895802
Rh001_022_010-    i_022    tia_h_in_001_010-    120572.06091277403
Rh001_023_010+    i_023    tia_h_in_001_010+    5000
Rh001_023_010-    i_023    tia_h_in_001_010-    53481.367851003786
Rh001_024_010+    i_024    tia_h_in_001_010+    119257.29177781288
Rh001_024_010-    i_024    tia_h_in_001_010-    78802.71758159524
Rh001_025_010+    i_025    tia_h_in_001_010+    121495.95010856965
Rh001_025_010-    i_025    tia_h_in_001_010-    91641.83046725592
Rh001_026_010+    i_026    tia_h_in_001_010+    121041.03692451582
Rh001_026_010-    i_026    tia_h_in_001_010-    56901.15838859207
Rh001_027_010+    i_027    tia_h_in_001_010+    5000
Rh001_027_010-    i_027    tia_h_in_001_010-    64010.53329669906
Rh001_028_010+    i_028    tia_h_in_001_010+    5000
Rh001_028_010-    i_028    tia_h_in_001_010-    96553.18015488771
Rh001_029_010+    i_029    tia_h_in_001_010+    5000
Rh001_029_010-    i_029    tia_h_in_001_010-    120089.24477720866
Rh001_030_010+    i_030    tia_h_in_001_010+    55790.936875077874
Rh001_030_010-    i_030    tia_h_in_001_010-    120082.22794837841
Rh001_031_010+    i_031    tia_h_in_001_010+    120000
Rh001_031_010-    i_031    tia_h_in_001_010-    120273.63397025251
Rh001_032_010+    i_032    tia_h_in_001_010+    118980.23252931518
Rh001_032_010-    i_032    tia_h_in_001_010-    67202.00514725863
Rh001_033_010+    i_033    tia_h_in_001_010+    121568.87811543905
Rh001_033_010-    i_033    tia_h_in_001_010-    63574.03000775955
Rh001_034_010+    i_034    tia_h_in_001_010+    58614.02754536625
Rh001_034_010-    i_034    tia_h_in_001_010-    118966.12486571973
Rh001_035_010+    i_035    tia_h_in_001_010+    86471.44238029157
Rh001_035_010-    i_035    tia_h_in_001_010-    120901.72275727348
Rh001_036_010+    i_036    tia_h_in_001_010+    119843.7965403959
Rh001_036_010-    i_036    tia_h_in_001_010-    117960.2150601392
Rh001_037_010+    i_037    tia_h_in_001_010+    105443.59227845771
Rh001_037_010-    i_037    tia_h_in_001_010-    122138.31719970504
Rh001_038_010+    i_038    tia_h_in_001_010+    119839.74847741723
Rh001_038_010-    i_038    tia_h_in_001_010-    58942.56462663801
Rh001_039_010+    i_039    tia_h_in_001_010+    121298.49429432275
Rh001_039_010-    i_039    tia_h_in_001_010-    5000
Rh001_040_010+    i_040    tia_h_in_001_010+    56105.285774761905
Rh001_040_010-    i_040    tia_h_in_001_010-    120643.6194176992
Rh001_041_010+    i_041    tia_h_in_001_010+    120000
Rh001_041_010-    i_041    tia_h_in_001_010-    88570.9994569131
Rh001_042_010+    i_042    tia_h_in_001_010+    119401.89554577909
Rh001_042_010-    i_042    tia_h_in_001_010-    107784.53965737818
Rh001_043_010+    i_043    tia_h_in_001_010+    119508.22192444475
Rh001_043_010-    i_043    tia_h_in_001_010-    57981.61862122081
Rh001_044_010+    i_044    tia_h_in_001_010+    121812.55955664688
Rh001_044_010-    i_044    tia_h_in_001_010-    68853.17658228143
Rh001_045_010+    i_045    tia_h_in_001_010+    120629.67021283641
Rh001_045_010-    i_045    tia_h_in_001_010-    111645.21577862906
Rh001_046_010+    i_046    tia_h_in_001_010+    121134.83506289922
Rh001_046_010-    i_046    tia_h_in_001_010-    65404.91317560655
Rh001_047_010+    i_047    tia_h_in_001_010+    121660.55858977888
Rh001_047_010-    i_047    tia_h_in_001_010-    101099.23849144593
Rh001_048_010+    i_048    tia_h_in_001_010+    82086.07989336789
Rh001_048_010-    i_048    tia_h_in_001_010-    120334.95568510013
Rh001_049_010+    i_049    tia_h_in_001_010+    5000
Rh001_049_010-    i_049    tia_h_in_001_010-    53127.650101829764
Rh001_050_010+    i_050    tia_h_in_001_010+    91440.66178141843
Rh001_050_010-    i_050    tia_h_in_001_010-    120309.82664798164
Rh001_051_010+    i_051    tia_h_in_001_010+    118711.61412293
Rh001_051_010-    i_051    tia_h_in_001_010-    64630.17152574909
Rh001_052_010+    i_052    tia_h_in_001_010+    121160.32252580307
Rh001_052_010-    i_052    tia_h_in_001_010-    73270.21637266631
Rh001_053_010+    i_053    tia_h_in_001_010+    120000
Rh001_053_010-    i_053    tia_h_in_001_010-    118905.02488382727
Rh001_054_010+    i_054    tia_h_in_001_010+    61341.52827042915
Rh001_054_010-    i_054    tia_h_in_001_010-    5000
Rh001_055_010+    i_055    tia_h_in_001_010+    120886.1808703955
Rh001_055_010-    i_055    tia_h_in_001_010-    84699.62173013562
Rh001_056_010+    i_056    tia_h_in_001_010+    118966.09319502328
Rh001_056_010-    i_056    tia_h_in_001_010-    76926.0068740911
Rh001_057_010+    i_057    tia_h_in_001_010+    119596.80485269663
Rh001_057_010-    i_057    tia_h_in_001_010-    55421.276189483666
Rh001_058_010+    i_058    tia_h_in_001_010+    5000
Rh001_058_010-    i_058    tia_h_in_001_010-    5000
Rh001_059_010+    i_059    tia_h_in_001_010+    119437.881565264
Rh001_059_010-    i_059    tia_h_in_001_010-    56478.23397223871
Rh001_060_010+    i_060    tia_h_in_001_010+    121210.6281650641
Rh001_060_010-    i_060    tia_h_in_001_010-    90238.63917431467
Rh001_061_010+    i_061    tia_h_in_001_010+    100260.42247425372
Rh001_061_010-    i_061    tia_h_in_001_010-    119911.11748579853
Rh001_062_010+    i_062    tia_h_in_001_010+    121960.21428707693
Rh001_062_010-    i_062    tia_h_in_001_010-    54112.29881014219
Rh001_063_010+    i_063    tia_h_in_001_010+    58204.87466018117
Rh001_063_010-    i_063    tia_h_in_001_010-    120324.97738831706
Rh001_064_010+    i_064    tia_h_in_001_010+    69565.33098416906
Rh001_064_010-    i_064    tia_h_in_001_010-    122701.10419372364

* Neuron 11
Rh001_001_011+    i_001    tia_h_in_001_011+    119552.54442684262
Rh001_001_011-    i_001    tia_h_in_001_011-    15093.855922997893
Rh001_002_011+    i_002    tia_h_in_001_011+    121164.69173840737
Rh001_002_011-    i_002    tia_h_in_001_011-    27595.985911656986
Rh001_003_011+    i_003    tia_h_in_001_011+    121255.01320280186
Rh001_003_011-    i_003    tia_h_in_001_011-    29954.511029647227
Rh001_004_011+    i_004    tia_h_in_001_011+    118367.16058883678
Rh001_004_011-    i_004    tia_h_in_001_011-    27002.243834645687
Rh001_005_011+    i_005    tia_h_in_001_011+    118376.93980814965
Rh001_005_011-    i_005    tia_h_in_001_011-    35488.82927327659
Rh001_006_011+    i_006    tia_h_in_001_011+    120082.35622124332
Rh001_006_011-    i_006    tia_h_in_001_011-    29111.255735993673
Rh001_007_011+    i_007    tia_h_in_001_011+    81939.90755749607
Rh001_007_011-    i_007    tia_h_in_001_011-    5000
Rh001_008_011+    i_008    tia_h_in_001_011+    119247.881391973
Rh001_008_011-    i_008    tia_h_in_001_011-    107026.42276744092
Rh001_009_011+    i_009    tia_h_in_001_011+    39258.98422440426
Rh001_009_011-    i_009    tia_h_in_001_011-    118943.56366970937
Rh001_010_011+    i_010    tia_h_in_001_011+    40536.418330698725
Rh001_010_011-    i_010    tia_h_in_001_011-    119564.00152984937
Rh001_011_011+    i_011    tia_h_in_001_011+    120000
Rh001_011_011-    i_011    tia_h_in_001_011-    120343.33954590232
Rh001_012_011+    i_012    tia_h_in_001_011+    33786.28121326111
Rh001_012_011-    i_012    tia_h_in_001_011-    120220.4680414818
Rh001_013_011+    i_013    tia_h_in_001_011+    72218.84705998408
Rh001_013_011-    i_013    tia_h_in_001_011-    117936.68087866476
Rh001_014_011+    i_014    tia_h_in_001_011+    122600.05282636927
Rh001_014_011-    i_014    tia_h_in_001_011-    97258.28732336909
Rh001_015_011+    i_015    tia_h_in_001_011+    120445.82374824719
Rh001_015_011-    i_015    tia_h_in_001_011-    55483.015307991336
Rh001_016_011+    i_016    tia_h_in_001_011+    120000
Rh001_016_011-    i_016    tia_h_in_001_011-    72703.214771108
Rh001_017_011+    i_017    tia_h_in_001_011+    39531.55188147452
Rh001_017_011-    i_017    tia_h_in_001_011-    119110.84867132032
Rh001_018_011+    i_018    tia_h_in_001_011+    37077.66341892743
Rh001_018_011-    i_018    tia_h_in_001_011-    121475.52366208786
Rh001_019_011+    i_019    tia_h_in_001_011+    121159.73370201654
Rh001_019_011-    i_019    tia_h_in_001_011-    57702.344904786645
Rh001_020_011+    i_020    tia_h_in_001_011+    43988.801440810435
Rh001_020_011-    i_020    tia_h_in_001_011-    118351.44125190031
Rh001_021_011+    i_021    tia_h_in_001_011+    27105.93077446599
Rh001_021_011-    i_021    tia_h_in_001_011-    120693.9372634427
Rh001_022_011+    i_022    tia_h_in_001_011+    73243.41555717244
Rh001_022_011-    i_022    tia_h_in_001_011-    120929.86997484976
Rh001_023_011+    i_023    tia_h_in_001_011+    119412.09464027476
Rh001_023_011-    i_023    tia_h_in_001_011-    115844.3054890412
Rh001_024_011+    i_024    tia_h_in_001_011+    86505.8651750201
Rh001_024_011-    i_024    tia_h_in_001_011-    117565.29634676824
Rh001_025_011+    i_025    tia_h_in_001_011+    52851.925503166894
Rh001_025_011-    i_025    tia_h_in_001_011-    120000
Rh001_026_011+    i_026    tia_h_in_001_011+    120145.58695098726
Rh001_026_011-    i_026    tia_h_in_001_011-    120000
Rh001_027_011+    i_027    tia_h_in_001_011+    120000
Rh001_027_011-    i_027    tia_h_in_001_011-    109288.75404452198
Rh001_028_011+    i_028    tia_h_in_001_011+    73152.62119123866
Rh001_028_011-    i_028    tia_h_in_001_011-    120406.37328827954
Rh001_029_011+    i_029    tia_h_in_001_011+    85685.55692993701
Rh001_029_011-    i_029    tia_h_in_001_011-    120349.53985238486
Rh001_030_011+    i_030    tia_h_in_001_011+    69383.3732416168
Rh001_030_011-    i_030    tia_h_in_001_011-    120888.94381704748
Rh001_031_011+    i_031    tia_h_in_001_011+    50489.85859575251
Rh001_031_011-    i_031    tia_h_in_001_011-    120033.93121079326
Rh001_032_011+    i_032    tia_h_in_001_011+    71877.25848055817
Rh001_032_011-    i_032    tia_h_in_001_011-    5000
Rh001_033_011+    i_033    tia_h_in_001_011+    120058.41176402502
Rh001_033_011-    i_033    tia_h_in_001_011-    96521.36220829892
Rh001_034_011+    i_034    tia_h_in_001_011+    120000
Rh001_034_011-    i_034    tia_h_in_001_011-    119417.78305988136
Rh001_035_011+    i_035    tia_h_in_001_011+    5000
Rh001_035_011-    i_035    tia_h_in_001_011-    119331.07016157283
Rh001_036_011+    i_036    tia_h_in_001_011+    119767.03450924144
Rh001_036_011-    i_036    tia_h_in_001_011-    32399.654014650718
Rh001_037_011+    i_037    tia_h_in_001_011+    121105.3011028137
Rh001_037_011-    i_037    tia_h_in_001_011-    104884.96957511538
Rh001_038_011+    i_038    tia_h_in_001_011+    57623.047086773106
Rh001_038_011-    i_038    tia_h_in_001_011-    5000
Rh001_039_011+    i_039    tia_h_in_001_011+    57433.53940782515
Rh001_039_011-    i_039    tia_h_in_001_011-    119839.85313289647
Rh001_040_011+    i_040    tia_h_in_001_011+    120000
Rh001_040_011-    i_040    tia_h_in_001_011-    38178.58516994328
Rh001_041_011+    i_041    tia_h_in_001_011+    77671.75991108827
Rh001_041_011-    i_041    tia_h_in_001_011-    119316.01711970972
Rh001_042_011+    i_042    tia_h_in_001_011+    120514.13683906106
Rh001_042_011-    i_042    tia_h_in_001_011-    117950.81106724226
Rh001_043_011+    i_043    tia_h_in_001_011+    120927.06367251895
Rh001_043_011-    i_043    tia_h_in_001_011-    44164.03240777733
Rh001_044_011+    i_044    tia_h_in_001_011+    119391.1256872149
Rh001_044_011-    i_044    tia_h_in_001_011-    51136.21849624475
Rh001_045_011+    i_045    tia_h_in_001_011+    119120.49939682214
Rh001_045_011-    i_045    tia_h_in_001_011-    34467.914090538114
Rh001_046_011+    i_046    tia_h_in_001_011+    120064.12498738634
Rh001_046_011-    i_046    tia_h_in_001_011-    50851.09399889871
Rh001_047_011+    i_047    tia_h_in_001_011+    58907.82375278527
Rh001_047_011-    i_047    tia_h_in_001_011-    119783.82509390028
Rh001_048_011+    i_048    tia_h_in_001_011+    119596.58777782504
Rh001_048_011-    i_048    tia_h_in_001_011-    5000
Rh001_049_011+    i_049    tia_h_in_001_011+    119698.89045469492
Rh001_049_011-    i_049    tia_h_in_001_011-    62651.33556469114
Rh001_050_011+    i_050    tia_h_in_001_011+    71474.91306784318
Rh001_050_011-    i_050    tia_h_in_001_011-    120549.54631434186
Rh001_051_011+    i_051    tia_h_in_001_011+    70616.27305829126
Rh001_051_011-    i_051    tia_h_in_001_011-    120419.04311963276
Rh001_052_011+    i_052    tia_h_in_001_011+    120000
Rh001_052_011-    i_052    tia_h_in_001_011-    121646.68779960032
Rh001_053_011+    i_053    tia_h_in_001_011+    54482.94456944134
Rh001_053_011-    i_053    tia_h_in_001_011-    117870.7732457774
Rh001_054_011+    i_054    tia_h_in_001_011+    5000
Rh001_054_011-    i_054    tia_h_in_001_011-    79836.33998756405
Rh001_055_011+    i_055    tia_h_in_001_011+    119243.12808861746
Rh001_055_011-    i_055    tia_h_in_001_011-    34536.66967630469
Rh001_056_011+    i_056    tia_h_in_001_011+    62168.1924305716
Rh001_056_011-    i_056    tia_h_in_001_011-    119572.5733553352
Rh001_057_011+    i_057    tia_h_in_001_011+    79894.71760884777
Rh001_057_011-    i_057    tia_h_in_001_011-    118660.63284384726
Rh001_058_011+    i_058    tia_h_in_001_011+    119471.24333105287
Rh001_058_011-    i_058    tia_h_in_001_011-    86774.2101222199
Rh001_059_011+    i_059    tia_h_in_001_011+    47330.40010110505
Rh001_059_011-    i_059    tia_h_in_001_011-    118838.37488529462
Rh001_060_011+    i_060    tia_h_in_001_011+    119586.92291792537
Rh001_060_011-    i_060    tia_h_in_001_011-    118295.19624253984
Rh001_061_011+    i_061    tia_h_in_001_011+    72324.0380148896
Rh001_061_011-    i_061    tia_h_in_001_011-    119505.04126019444
Rh001_062_011+    i_062    tia_h_in_001_011+    118604.7869652056
Rh001_062_011-    i_062    tia_h_in_001_011-    87828.88830614119
Rh001_063_011+    i_063    tia_h_in_001_011+    39315.66413689932
Rh001_063_011-    i_063    tia_h_in_001_011-    120750.24719407078
Rh001_064_011+    i_064    tia_h_in_001_011+    120622.05135904693
Rh001_064_011-    i_064    tia_h_in_001_011-    96204.01016672322

* Neuron 12
Rh001_001_012+    i_001    tia_h_in_001_012+    120390.35994256036
Rh001_001_012-    i_001    tia_h_in_001_012-    29728.23085890002
Rh001_002_012+    i_002    tia_h_in_001_012+    120000
Rh001_002_012-    i_002    tia_h_in_001_012-    120000
Rh001_003_012+    i_003    tia_h_in_001_012+    5000
Rh001_003_012-    i_003    tia_h_in_001_012-    30423.098726773813
Rh001_004_012+    i_004    tia_h_in_001_012+    120000
Rh001_004_012-    i_004    tia_h_in_001_012-    5000
Rh001_005_012+    i_005    tia_h_in_001_012+    59747.813011295635
Rh001_005_012-    i_005    tia_h_in_001_012-    120675.63182055455
Rh001_006_012+    i_006    tia_h_in_001_012+    120000
Rh001_006_012-    i_006    tia_h_in_001_012-    51577.28781015271
Rh001_007_012+    i_007    tia_h_in_001_012+    117353.96826405032
Rh001_007_012-    i_007    tia_h_in_001_012-    119756.08567812179
Rh001_008_012+    i_008    tia_h_in_001_012+    120000
Rh001_008_012-    i_008    tia_h_in_001_012-    93752.3002614206
Rh001_009_012+    i_009    tia_h_in_001_012+    92441.1259587011
Rh001_009_012-    i_009    tia_h_in_001_012-    5000
Rh001_010_012+    i_010    tia_h_in_001_012+    5000
Rh001_010_012-    i_010    tia_h_in_001_012-    32774.77236131687
Rh001_011_012+    i_011    tia_h_in_001_012+    120266.59715513002
Rh001_011_012-    i_011    tia_h_in_001_012-    58428.71899380737
Rh001_012_012+    i_012    tia_h_in_001_012+    121788.97420553467
Rh001_012_012-    i_012    tia_h_in_001_012-    36426.836774662
Rh001_013_012+    i_013    tia_h_in_001_012+    5000
Rh001_013_012-    i_013    tia_h_in_001_012-    119941.97826526704
Rh001_014_012+    i_014    tia_h_in_001_012+    41978.92603694759
Rh001_014_012-    i_014    tia_h_in_001_012-    119132.04466511584
Rh001_015_012+    i_015    tia_h_in_001_012+    68773.42669299609
Rh001_015_012-    i_015    tia_h_in_001_012-    119158.80553785774
Rh001_016_012+    i_016    tia_h_in_001_012+    91797.420328266
Rh001_016_012-    i_016    tia_h_in_001_012-    118854.39160545164
Rh001_017_012+    i_017    tia_h_in_001_012+    120671.60768538789
Rh001_017_012-    i_017    tia_h_in_001_012-    53282.09307053081
Rh001_018_012+    i_018    tia_h_in_001_012+    39254.70836589518
Rh001_018_012-    i_018    tia_h_in_001_012-    120000
Rh001_019_012+    i_019    tia_h_in_001_012+    80307.09333266104
Rh001_019_012-    i_019    tia_h_in_001_012-    119244.40416246897
Rh001_020_012+    i_020    tia_h_in_001_012+    119746.82677980266
Rh001_020_012-    i_020    tia_h_in_001_012-    26118.9232443771
Rh001_021_012+    i_021    tia_h_in_001_012+    119587.03070744242
Rh001_021_012-    i_021    tia_h_in_001_012-    85807.02011343351
Rh001_022_012+    i_022    tia_h_in_001_012+    121011.35923943503
Rh001_022_012-    i_022    tia_h_in_001_012-    52787.07913625172
Rh001_023_012+    i_023    tia_h_in_001_012+    40853.48423530765
Rh001_023_012-    i_023    tia_h_in_001_012-    120628.15932405234
Rh001_024_012+    i_024    tia_h_in_001_012+    119422.62012513082
Rh001_024_012-    i_024    tia_h_in_001_012-    79398.28519443305
Rh001_025_012+    i_025    tia_h_in_001_012+    120405.26841805634
Rh001_025_012-    i_025    tia_h_in_001_012-    37628.32973057253
Rh001_026_012+    i_026    tia_h_in_001_012+    82873.12473591862
Rh001_026_012-    i_026    tia_h_in_001_012-    121937.18978988353
Rh001_027_012+    i_027    tia_h_in_001_012+    38230.18479769309
Rh001_027_012-    i_027    tia_h_in_001_012-    121382.74064694889
Rh001_028_012+    i_028    tia_h_in_001_012+    56422.579525524656
Rh001_028_012-    i_028    tia_h_in_001_012-    119582.1785534281
Rh001_029_012+    i_029    tia_h_in_001_012+    121194.17407672184
Rh001_029_012-    i_029    tia_h_in_001_012-    83215.7395404768
Rh001_030_012+    i_030    tia_h_in_001_012+    120000
Rh001_030_012-    i_030    tia_h_in_001_012-    77932.16059797916
Rh001_031_012+    i_031    tia_h_in_001_012+    43274.86396562979
Rh001_031_012-    i_031    tia_h_in_001_012-    121240.44087616623
Rh001_032_012+    i_032    tia_h_in_001_012+    26494.41007274848
Rh001_032_012-    i_032    tia_h_in_001_012-    119811.81881484973
Rh001_033_012+    i_033    tia_h_in_001_012+    43579.83162786385
Rh001_033_012-    i_033    tia_h_in_001_012-    120067.14874632814
Rh001_034_012+    i_034    tia_h_in_001_012+    120704.20449611139
Rh001_034_012-    i_034    tia_h_in_001_012-    112125.94746517684
Rh001_035_012+    i_035    tia_h_in_001_012+    58216.99249374424
Rh001_035_012-    i_035    tia_h_in_001_012-    120128.30595519004
Rh001_036_012+    i_036    tia_h_in_001_012+    120000
Rh001_036_012-    i_036    tia_h_in_001_012-    120398.09623127646
Rh001_037_012+    i_037    tia_h_in_001_012+    120000
Rh001_037_012-    i_037    tia_h_in_001_012-    119312.51814295736
Rh001_038_012+    i_038    tia_h_in_001_012+    92768.61511009473
Rh001_038_012-    i_038    tia_h_in_001_012-    120468.93893054096
Rh001_039_012+    i_039    tia_h_in_001_012+    63212.75739314751
Rh001_039_012-    i_039    tia_h_in_001_012-    121671.72178397125
Rh001_040_012+    i_040    tia_h_in_001_012+    119766.76565093317
Rh001_040_012-    i_040    tia_h_in_001_012-    50938.25759817771
Rh001_041_012+    i_041    tia_h_in_001_012+    35591.8624484636
Rh001_041_012-    i_041    tia_h_in_001_012-    121002.86421047719
Rh001_042_012+    i_042    tia_h_in_001_012+    57849.89978881952
Rh001_042_012-    i_042    tia_h_in_001_012-    119240.37500357792
Rh001_043_012+    i_043    tia_h_in_001_012+    114070.34073960557
Rh001_043_012-    i_043    tia_h_in_001_012-    120477.41483533313
Rh001_044_012+    i_044    tia_h_in_001_012+    120000
Rh001_044_012-    i_044    tia_h_in_001_012-    121497.82445407577
Rh001_045_012+    i_045    tia_h_in_001_012+    119378.39864703687
Rh001_045_012-    i_045    tia_h_in_001_012-    47649.92639711713
Rh001_046_012+    i_046    tia_h_in_001_012+    5000
Rh001_046_012-    i_046    tia_h_in_001_012-    42384.03297940924
Rh001_047_012+    i_047    tia_h_in_001_012+    74125.54314156681
Rh001_047_012-    i_047    tia_h_in_001_012-    119335.69517172973
Rh001_048_012+    i_048    tia_h_in_001_012+    120978.4945510349
Rh001_048_012-    i_048    tia_h_in_001_012-    40895.639890423794
Rh001_049_012+    i_049    tia_h_in_001_012+    42470.156239439435
Rh001_049_012-    i_049    tia_h_in_001_012-    121252.22727955303
Rh001_050_012+    i_050    tia_h_in_001_012+    120000
Rh001_050_012-    i_050    tia_h_in_001_012-    120000
Rh001_051_012+    i_051    tia_h_in_001_012+    120114.85846205954
Rh001_051_012-    i_051    tia_h_in_001_012-    79829.15893350846
Rh001_052_012+    i_052    tia_h_in_001_012+    79772.53879490077
Rh001_052_012-    i_052    tia_h_in_001_012-    120148.86507983667
Rh001_053_012+    i_053    tia_h_in_001_012+    5000
Rh001_053_012-    i_053    tia_h_in_001_012-    119344.4186048379
Rh001_054_012+    i_054    tia_h_in_001_012+    66345.73654436994
Rh001_054_012-    i_054    tia_h_in_001_012-    121539.74698254955
Rh001_055_012+    i_055    tia_h_in_001_012+    120000
Rh001_055_012-    i_055    tia_h_in_001_012-    45393.3530695167
Rh001_056_012+    i_056    tia_h_in_001_012+    117250.84138220956
Rh001_056_012-    i_056    tia_h_in_001_012-    120357.60526435198
Rh001_057_012+    i_057    tia_h_in_001_012+    119111.4249593581
Rh001_057_012-    i_057    tia_h_in_001_012-    44225.36004525714
Rh001_058_012+    i_058    tia_h_in_001_012+    89961.70687891521
Rh001_058_012-    i_058    tia_h_in_001_012-    120768.03384585495
Rh001_059_012+    i_059    tia_h_in_001_012+    120068.40587248381
Rh001_059_012-    i_059    tia_h_in_001_012-    49493.90202988661
Rh001_060_012+    i_060    tia_h_in_001_012+    120339.12710132859
Rh001_060_012-    i_060    tia_h_in_001_012-    46598.848570586575
Rh001_061_012+    i_061    tia_h_in_001_012+    66778.00167511123
Rh001_061_012-    i_061    tia_h_in_001_012-    121069.3040283728
Rh001_062_012+    i_062    tia_h_in_001_012+    120000
Rh001_062_012-    i_062    tia_h_in_001_012-    42000.49588367603
Rh001_063_012+    i_063    tia_h_in_001_012+    120724.00524975474
Rh001_063_012-    i_063    tia_h_in_001_012-    120000
Rh001_064_012+    i_064    tia_h_in_001_012+    121495.09024036366
Rh001_064_012-    i_064    tia_h_in_001_012-    58828.1528860639

* Neuron 13
Rh001_001_013+    i_001    tia_h_in_001_013+    120692.4251947382
Rh001_001_013-    i_001    tia_h_in_001_013-    5000
Rh001_002_013+    i_002    tia_h_in_001_013+    121580.5754208126
Rh001_002_013-    i_002    tia_h_in_001_013-    16812.052604756384
Rh001_003_013+    i_003    tia_h_in_001_013+    120819.91108005881
Rh001_003_013-    i_003    tia_h_in_001_013-    33735.49443828539
Rh001_004_013+    i_004    tia_h_in_001_013+    121030.24281565452
Rh001_004_013-    i_004    tia_h_in_001_013-    36721.41109695026
Rh001_005_013+    i_005    tia_h_in_001_013+    121239.979133596
Rh001_005_013-    i_005    tia_h_in_001_013-    5000
Rh001_006_013+    i_006    tia_h_in_001_013+    52001.37531470694
Rh001_006_013-    i_006    tia_h_in_001_013-    5000
Rh001_007_013+    i_007    tia_h_in_001_013+    5000
Rh001_007_013-    i_007    tia_h_in_001_013-    61394.32805023102
Rh001_008_013+    i_008    tia_h_in_001_013+    57601.35728098991
Rh001_008_013-    i_008    tia_h_in_001_013-    120701.39871524795
Rh001_009_013+    i_009    tia_h_in_001_013+    71583.580733036
Rh001_009_013-    i_009    tia_h_in_001_013-    118787.73040846887
Rh001_010_013+    i_010    tia_h_in_001_013+    120000
Rh001_010_013-    i_010    tia_h_in_001_013-    120818.2323557111
Rh001_011_013+    i_011    tia_h_in_001_013+    43427.17909271055
Rh001_011_013-    i_011    tia_h_in_001_013-    119159.96856686818
Rh001_012_013+    i_012    tia_h_in_001_013+    120492.45023750076
Rh001_012_013-    i_012    tia_h_in_001_013-    58474.69391991533
Rh001_013_013+    i_013    tia_h_in_001_013+    5000
Rh001_013_013-    i_013    tia_h_in_001_013-    101812.97049396978
Rh001_014_013+    i_014    tia_h_in_001_013+    119679.63423492374
Rh001_014_013-    i_014    tia_h_in_001_013-    56512.71753355149
Rh001_015_013+    i_015    tia_h_in_001_013+    92585.17696319474
Rh001_015_013-    i_015    tia_h_in_001_013-    120762.71219469771
Rh001_016_013+    i_016    tia_h_in_001_013+    77451.17668820477
Rh001_016_013-    i_016    tia_h_in_001_013-    118906.61723041031
Rh001_017_013+    i_017    tia_h_in_001_013+    21864.276415924232
Rh001_017_013-    i_017    tia_h_in_001_013-    119700.76098294473
Rh001_018_013+    i_018    tia_h_in_001_013+    36874.23035955973
Rh001_018_013-    i_018    tia_h_in_001_013-    120357.68382475973
Rh001_019_013+    i_019    tia_h_in_001_013+    40952.690063295464
Rh001_019_013-    i_019    tia_h_in_001_013-    121414.8912408357
Rh001_020_013+    i_020    tia_h_in_001_013+    97570.37870558209
Rh001_020_013-    i_020    tia_h_in_001_013-    120374.57197355911
Rh001_021_013+    i_021    tia_h_in_001_013+    117828.58184062886
Rh001_021_013-    i_021    tia_h_in_001_013-    67234.65278340412
Rh001_022_013+    i_022    tia_h_in_001_013+    118497.81686886276
Rh001_022_013-    i_022    tia_h_in_001_013-    59784.204777276944
Rh001_023_013+    i_023    tia_h_in_001_013+    119553.27844922832
Rh001_023_013-    i_023    tia_h_in_001_013-    45575.2989466466
Rh001_024_013+    i_024    tia_h_in_001_013+    120322.14559846757
Rh001_024_013-    i_024    tia_h_in_001_013-    29175.28407152177
Rh001_025_013+    i_025    tia_h_in_001_013+    5000
Rh001_025_013-    i_025    tia_h_in_001_013-    119611.18855457782
Rh001_026_013+    i_026    tia_h_in_001_013+    63963.824316393984
Rh001_026_013-    i_026    tia_h_in_001_013-    120646.36970770858
Rh001_027_013+    i_027    tia_h_in_001_013+    51164.93288162605
Rh001_027_013-    i_027    tia_h_in_001_013-    119469.7577831696
Rh001_028_013+    i_028    tia_h_in_001_013+    120000
Rh001_028_013-    i_028    tia_h_in_001_013-    5000
Rh001_029_013+    i_029    tia_h_in_001_013+    119277.65907357693
Rh001_029_013-    i_029    tia_h_in_001_013-    34479.229591897725
Rh001_030_013+    i_030    tia_h_in_001_013+    63808.100964034544
Rh001_030_013-    i_030    tia_h_in_001_013-    5000
Rh001_031_013+    i_031    tia_h_in_001_013+    119434.71564455878
Rh001_031_013-    i_031    tia_h_in_001_013-    74510.5535631733
Rh001_032_013+    i_032    tia_h_in_001_013+    67707.30603113842
Rh001_032_013-    i_032    tia_h_in_001_013-    119898.79743662204
Rh001_033_013+    i_033    tia_h_in_001_013+    5000
Rh001_033_013-    i_033    tia_h_in_001_013-    72288.13580666836
Rh001_034_013+    i_034    tia_h_in_001_013+    120209.61390664199
Rh001_034_013-    i_034    tia_h_in_001_013-    62819.73617820218
Rh001_035_013+    i_035    tia_h_in_001_013+    120193.41168647645
Rh001_035_013-    i_035    tia_h_in_001_013-    97108.38137761071
Rh001_036_013+    i_036    tia_h_in_001_013+    5000
Rh001_036_013-    i_036    tia_h_in_001_013-    5000
Rh001_037_013+    i_037    tia_h_in_001_013+    33226.841155269336
Rh001_037_013-    i_037    tia_h_in_001_013-    118990.29385012061
Rh001_038_013+    i_038    tia_h_in_001_013+    5000
Rh001_038_013-    i_038    tia_h_in_001_013-    120000
Rh001_039_013+    i_039    tia_h_in_001_013+    120000
Rh001_039_013-    i_039    tia_h_in_001_013-    120909.88621849888
Rh001_040_013+    i_040    tia_h_in_001_013+    121031.83589767902
Rh001_040_013-    i_040    tia_h_in_001_013-    59746.6139511552
Rh001_041_013+    i_041    tia_h_in_001_013+    121317.2205060229
Rh001_041_013-    i_041    tia_h_in_001_013-    63109.118990103234
Rh001_042_013+    i_042    tia_h_in_001_013+    79075.43512255138
Rh001_042_013-    i_042    tia_h_in_001_013-    118919.56129140593
Rh001_043_013+    i_043    tia_h_in_001_013+    116007.16473182123
Rh001_043_013-    i_043    tia_h_in_001_013-    120921.63703046052
Rh001_044_013+    i_044    tia_h_in_001_013+    101296.1806107937
Rh001_044_013-    i_044    tia_h_in_001_013-    119732.8676779085
Rh001_045_013+    i_045    tia_h_in_001_013+    29760.07350244263
Rh001_045_013-    i_045    tia_h_in_001_013-    121577.13375130802
Rh001_046_013+    i_046    tia_h_in_001_013+    33410.959645607014
Rh001_046_013-    i_046    tia_h_in_001_013-    120000
Rh001_047_013+    i_047    tia_h_in_001_013+    120000
Rh001_047_013-    i_047    tia_h_in_001_013-    119150.94578109389
Rh001_048_013+    i_048    tia_h_in_001_013+    118279.24721398026
Rh001_048_013-    i_048    tia_h_in_001_013-    84129.01752535213
Rh001_049_013+    i_049    tia_h_in_001_013+    119845.30128113637
Rh001_049_013-    i_049    tia_h_in_001_013-    64855.07154236718
Rh001_050_013+    i_050    tia_h_in_001_013+    119695.10034146636
Rh001_050_013-    i_050    tia_h_in_001_013-    98858.47578798574
Rh001_051_013+    i_051    tia_h_in_001_013+    98963.31215737022
Rh001_051_013-    i_051    tia_h_in_001_013-    121086.34059053307
Rh001_052_013+    i_052    tia_h_in_001_013+    118207.90303989605
Rh001_052_013-    i_052    tia_h_in_001_013-    57112.44713487979
Rh001_053_013+    i_053    tia_h_in_001_013+    118692.26117460089
Rh001_053_013-    i_053    tia_h_in_001_013-    59603.18155050884
Rh001_054_013+    i_054    tia_h_in_001_013+    56077.08819913569
Rh001_054_013-    i_054    tia_h_in_001_013-    118966.30892048219
Rh001_055_013+    i_055    tia_h_in_001_013+    69261.97483045387
Rh001_055_013-    i_055    tia_h_in_001_013-    120204.41356060424
Rh001_056_013+    i_056    tia_h_in_001_013+    93551.34915139708
Rh001_056_013-    i_056    tia_h_in_001_013-    120788.47196439755
Rh001_057_013+    i_057    tia_h_in_001_013+    120000
Rh001_057_013-    i_057    tia_h_in_001_013-    119483.11248123828
Rh001_058_013+    i_058    tia_h_in_001_013+    119795.7914689879
Rh001_058_013-    i_058    tia_h_in_001_013-    76372.00788617661
Rh001_059_013+    i_059    tia_h_in_001_013+    119140.97882445644
Rh001_059_013-    i_059    tia_h_in_001_013-    81045.3804374902
Rh001_060_013+    i_060    tia_h_in_001_013+    120000
Rh001_060_013-    i_060    tia_h_in_001_013-    121562.16796262535
Rh001_061_013+    i_061    tia_h_in_001_013+    119531.74721219219
Rh001_061_013-    i_061    tia_h_in_001_013-    99857.91423604253
Rh001_062_013+    i_062    tia_h_in_001_013+    118374.29398798819
Rh001_062_013-    i_062    tia_h_in_001_013-    76116.61868498744
Rh001_063_013+    i_063    tia_h_in_001_013+    120518.51057934522
Rh001_063_013-    i_063    tia_h_in_001_013-    46836.787093285464
Rh001_064_013+    i_064    tia_h_in_001_013+    50453.7841922504
Rh001_064_013-    i_064    tia_h_in_001_013-    120000

* Neuron 14
Rh001_001_014+    i_001    tia_h_in_001_014+    120657.41279524939
Rh001_001_014-    i_001    tia_h_in_001_014-    57340.17200372296
Rh001_002_014+    i_002    tia_h_in_001_014+    120369.52679412623
Rh001_002_014-    i_002    tia_h_in_001_014-    90946.33322050275
Rh001_003_014+    i_003    tia_h_in_001_014+    114261.81782462118
Rh001_003_014-    i_003    tia_h_in_001_014-    119416.65670443575
Rh001_004_014+    i_004    tia_h_in_001_014+    119616.85811265444
Rh001_004_014-    i_004    tia_h_in_001_014-    65160.16329164942
Rh001_005_014+    i_005    tia_h_in_001_014+    5000
Rh001_005_014-    i_005    tia_h_in_001_014-    120680.8494046178
Rh001_006_014+    i_006    tia_h_in_001_014+    118787.85662927416
Rh001_006_014-    i_006    tia_h_in_001_014-    48201.041972343024
Rh001_007_014+    i_007    tia_h_in_001_014+    120807.17682640062
Rh001_007_014-    i_007    tia_h_in_001_014-    56937.03002540676
Rh001_008_014+    i_008    tia_h_in_001_014+    5000
Rh001_008_014-    i_008    tia_h_in_001_014-    49913.414002270845
Rh001_009_014+    i_009    tia_h_in_001_014+    120374.34133925471
Rh001_009_014-    i_009    tia_h_in_001_014-    73879.20051636246
Rh001_010_014+    i_010    tia_h_in_001_014+    121538.67982567783
Rh001_010_014-    i_010    tia_h_in_001_014-    70151.38382686285
Rh001_011_014+    i_011    tia_h_in_001_014+    121240.45047216173
Rh001_011_014-    i_011    tia_h_in_001_014-    118770.55059357615
Rh001_012_014+    i_012    tia_h_in_001_014+    120174.79102017828
Rh001_012_014-    i_012    tia_h_in_001_014-    81434.03486330633
Rh001_013_014+    i_013    tia_h_in_001_014+    85149.23344759498
Rh001_013_014-    i_013    tia_h_in_001_014-    118674.09644519728
Rh001_014_014+    i_014    tia_h_in_001_014+    62157.0096338186
Rh001_014_014-    i_014    tia_h_in_001_014-    5000
Rh001_015_014+    i_015    tia_h_in_001_014+    99371.8142851751
Rh001_015_014-    i_015    tia_h_in_001_014-    118705.11179779157
Rh001_016_014+    i_016    tia_h_in_001_014+    117675.52106380386
Rh001_016_014-    i_016    tia_h_in_001_014-    65227.43686385339
Rh001_017_014+    i_017    tia_h_in_001_014+    120990.02487200062
Rh001_017_014-    i_017    tia_h_in_001_014-    52211.07962826887
Rh001_018_014+    i_018    tia_h_in_001_014+    92681.91827232209
Rh001_018_014-    i_018    tia_h_in_001_014-    120420.36707824147
Rh001_019_014+    i_019    tia_h_in_001_014+    119948.49395535637
Rh001_019_014-    i_019    tia_h_in_001_014-    68928.92798998626
Rh001_020_014+    i_020    tia_h_in_001_014+    5000
Rh001_020_014-    i_020    tia_h_in_001_014-    119647.55306266776
Rh001_021_014+    i_021    tia_h_in_001_014+    77481.54357253049
Rh001_021_014-    i_021    tia_h_in_001_014-    119153.9212568068
Rh001_022_014+    i_022    tia_h_in_001_014+    96213.90020668136
Rh001_022_014-    i_022    tia_h_in_001_014-    120287.91419313254
Rh001_023_014+    i_023    tia_h_in_001_014+    62494.351900639725
Rh001_023_014-    i_023    tia_h_in_001_014-    119002.04453938875
Rh001_024_014+    i_024    tia_h_in_001_014+    64097.18898062567
Rh001_024_014-    i_024    tia_h_in_001_014-    121555.90272160505
Rh001_025_014+    i_025    tia_h_in_001_014+    109450.44981620087
Rh001_025_014-    i_025    tia_h_in_001_014-    120717.05467022145
Rh001_026_014+    i_026    tia_h_in_001_014+    120865.5486825247
Rh001_026_014-    i_026    tia_h_in_001_014-    58594.95947725232
Rh001_027_014+    i_027    tia_h_in_001_014+    120000
Rh001_027_014-    i_027    tia_h_in_001_014-    121404.7130093057
Rh001_028_014+    i_028    tia_h_in_001_014+    118967.23773163628
Rh001_028_014-    i_028    tia_h_in_001_014-    120000
Rh001_029_014+    i_029    tia_h_in_001_014+    121048.87578634822
Rh001_029_014-    i_029    tia_h_in_001_014-    63201.72199140046
Rh001_030_014+    i_030    tia_h_in_001_014+    67027.10484502862
Rh001_030_014-    i_030    tia_h_in_001_014-    119938.67255353315
Rh001_031_014+    i_031    tia_h_in_001_014+    69356.34501476797
Rh001_031_014-    i_031    tia_h_in_001_014-    121180.43587281095
Rh001_032_014+    i_032    tia_h_in_001_014+    111788.06892650205
Rh001_032_014-    i_032    tia_h_in_001_014-    119524.09138381889
Rh001_033_014+    i_033    tia_h_in_001_014+    120110.37110954888
Rh001_033_014-    i_033    tia_h_in_001_014-    98138.34129915418
Rh001_034_014+    i_034    tia_h_in_001_014+    120268.47345211783
Rh001_034_014-    i_034    tia_h_in_001_014-    54877.858890082054
Rh001_035_014+    i_035    tia_h_in_001_014+    120195.90412933506
Rh001_035_014-    i_035    tia_h_in_001_014-    90703.21552267352
Rh001_036_014+    i_036    tia_h_in_001_014+    57343.85733981633
Rh001_036_014-    i_036    tia_h_in_001_014-    5000
Rh001_037_014+    i_037    tia_h_in_001_014+    111478.26226620746
Rh001_037_014-    i_037    tia_h_in_001_014-    119859.15216704519
Rh001_038_014+    i_038    tia_h_in_001_014+    120198.51544167336
Rh001_038_014-    i_038    tia_h_in_001_014-    107731.70124202092
Rh001_039_014+    i_039    tia_h_in_001_014+    5000
Rh001_039_014-    i_039    tia_h_in_001_014-    77956.66056087714
Rh001_040_014+    i_040    tia_h_in_001_014+    120385.47938953296
Rh001_040_014-    i_040    tia_h_in_001_014-    74266.07708496631
Rh001_041_014+    i_041    tia_h_in_001_014+    81470.51976183227
Rh001_041_014-    i_041    tia_h_in_001_014-    119878.73700617797
Rh001_042_014+    i_042    tia_h_in_001_014+    120543.59253331854
Rh001_042_014-    i_042    tia_h_in_001_014-    100023.42278883723
Rh001_043_014+    i_043    tia_h_in_001_014+    75953.4251201094
Rh001_043_014-    i_043    tia_h_in_001_014-    119856.44001805138
Rh001_044_014+    i_044    tia_h_in_001_014+    120532.95144089664
Rh001_044_014-    i_044    tia_h_in_001_014-    85987.42857448591
Rh001_045_014+    i_045    tia_h_in_001_014+    87970.38828721955
Rh001_045_014-    i_045    tia_h_in_001_014-    119747.7004299363
Rh001_046_014+    i_046    tia_h_in_001_014+    93393.74897108538
Rh001_046_014-    i_046    tia_h_in_001_014-    119826.01537894618
Rh001_047_014+    i_047    tia_h_in_001_014+    120718.16365442296
Rh001_047_014-    i_047    tia_h_in_001_014-    116280.30424111738
Rh001_048_014+    i_048    tia_h_in_001_014+    120000
Rh001_048_014-    i_048    tia_h_in_001_014-    120000
Rh001_049_014+    i_049    tia_h_in_001_014+    81779.56137497489
Rh001_049_014-    i_049    tia_h_in_001_014-    120338.94595502745
Rh001_050_014+    i_050    tia_h_in_001_014+    64821.57480096091
Rh001_050_014-    i_050    tia_h_in_001_014-    118344.10261097888
Rh001_051_014+    i_051    tia_h_in_001_014+    72682.40194044479
Rh001_051_014-    i_051    tia_h_in_001_014-    5000
Rh001_052_014+    i_052    tia_h_in_001_014+    119266.67369557987
Rh001_052_014-    i_052    tia_h_in_001_014-    74979.05365456502
Rh001_053_014+    i_053    tia_h_in_001_014+    120155.3179197779
Rh001_053_014-    i_053    tia_h_in_001_014-    52317.990925138816
Rh001_054_014+    i_054    tia_h_in_001_014+    5000
Rh001_054_014-    i_054    tia_h_in_001_014-    114495.91758753388
Rh001_055_014+    i_055    tia_h_in_001_014+    5000
Rh001_055_014-    i_055    tia_h_in_001_014-    98680.29526415559
Rh001_056_014+    i_056    tia_h_in_001_014+    119947.33339793707
Rh001_056_014-    i_056    tia_h_in_001_014-    82146.57602085035
Rh001_057_014+    i_057    tia_h_in_001_014+    120907.10952743526
Rh001_057_014-    i_057    tia_h_in_001_014-    77408.76543450446
Rh001_058_014+    i_058    tia_h_in_001_014+    121175.68922494343
Rh001_058_014-    i_058    tia_h_in_001_014-    92755.75826471986
Rh001_059_014+    i_059    tia_h_in_001_014+    74026.03378701802
Rh001_059_014-    i_059    tia_h_in_001_014-    119690.19248001746
Rh001_060_014+    i_060    tia_h_in_001_014+    111378.50604911518
Rh001_060_014-    i_060    tia_h_in_001_014-    121904.45199097968
Rh001_061_014+    i_061    tia_h_in_001_014+    120761.9973938202
Rh001_061_014-    i_061    tia_h_in_001_014-    72906.18983751649
Rh001_062_014+    i_062    tia_h_in_001_014+    120104.40538259404
Rh001_062_014-    i_062    tia_h_in_001_014-    68482.9874647947
Rh001_063_014+    i_063    tia_h_in_001_014+    119722.17118328647
Rh001_063_014-    i_063    tia_h_in_001_014-    82224.91691543347
Rh001_064_014+    i_064    tia_h_in_001_014+    119950.13997841832
Rh001_064_014-    i_064    tia_h_in_001_014-    70865.50924102713

* Neuron 15
Rh001_001_015+    i_001    tia_h_in_001_015+    58183.31841418034
Rh001_001_015-    i_001    tia_h_in_001_015-    5000
Rh001_002_015+    i_002    tia_h_in_001_015+    77501.7240352576
Rh001_002_015-    i_002    tia_h_in_001_015-    120017.34705674993
Rh001_003_015+    i_003    tia_h_in_001_015+    59377.68007521184
Rh001_003_015-    i_003    tia_h_in_001_015-    119252.71294018322
Rh001_004_015+    i_004    tia_h_in_001_015+    120356.27866286741
Rh001_004_015-    i_004    tia_h_in_001_015-    110073.42196924235
Rh001_005_015+    i_005    tia_h_in_001_015+    106062.66715872604
Rh001_005_015-    i_005    tia_h_in_001_015-    121559.13404884617
Rh001_006_015+    i_006    tia_h_in_001_015+    120000
Rh001_006_015-    i_006    tia_h_in_001_015-    119574.80409562714
Rh001_007_015+    i_007    tia_h_in_001_015+    119841.05513681985
Rh001_007_015-    i_007    tia_h_in_001_015-    52860.707775876945
Rh001_008_015+    i_008    tia_h_in_001_015+    120125.90419284676
Rh001_008_015-    i_008    tia_h_in_001_015-    119258.57551117026
Rh001_009_015+    i_009    tia_h_in_001_015+    119964.43452997661
Rh001_009_015-    i_009    tia_h_in_001_015-    102486.80320454459
Rh001_010_015+    i_010    tia_h_in_001_015+    120000
Rh001_010_015-    i_010    tia_h_in_001_015-    65579.40743806298
Rh001_011_015+    i_011    tia_h_in_001_015+    120220.17347996797
Rh001_011_015-    i_011    tia_h_in_001_015-    58117.56657752157
Rh001_012_015+    i_012    tia_h_in_001_015+    60276.50724085673
Rh001_012_015-    i_012    tia_h_in_001_015-    120377.0069284271
Rh001_013_015+    i_013    tia_h_in_001_015+    63059.62042255515
Rh001_013_015-    i_013    tia_h_in_001_015-    119005.89516150982
Rh001_014_015+    i_014    tia_h_in_001_015+    82520.32653653329
Rh001_014_015-    i_014    tia_h_in_001_015-    119428.8143951927
Rh001_015_015+    i_015    tia_h_in_001_015+    57716.39972597883
Rh001_015_015-    i_015    tia_h_in_001_015-    120207.51877760097
Rh001_016_015+    i_016    tia_h_in_001_015+    119556.54676346183
Rh001_016_015-    i_016    tia_h_in_001_015-    76082.39376087408
Rh001_017_015+    i_017    tia_h_in_001_015+    119716.53904914956
Rh001_017_015-    i_017    tia_h_in_001_015-    92578.62544643562
Rh001_018_015+    i_018    tia_h_in_001_015+    87898.27016355687
Rh001_018_015-    i_018    tia_h_in_001_015-    119274.67362056066
Rh001_019_015+    i_019    tia_h_in_001_015+    118670.12900043622
Rh001_019_015-    i_019    tia_h_in_001_015-    93696.09383990533
Rh001_020_015+    i_020    tia_h_in_001_015+    121178.50814855982
Rh001_020_015-    i_020    tia_h_in_001_015-    5000
Rh001_021_015+    i_021    tia_h_in_001_015+    5000
Rh001_021_015-    i_021    tia_h_in_001_015-    56366.306474920726
Rh001_022_015+    i_022    tia_h_in_001_015+    100263.30180037807
Rh001_022_015-    i_022    tia_h_in_001_015-    121083.38393955126
Rh001_023_015+    i_023    tia_h_in_001_015+    120283.13504432215
Rh001_023_015-    i_023    tia_h_in_001_015-    64504.264772137336
Rh001_024_015+    i_024    tia_h_in_001_015+    5000
Rh001_024_015-    i_024    tia_h_in_001_015-    116439.0841024915
Rh001_025_015+    i_025    tia_h_in_001_015+    56436.61372674748
Rh001_025_015-    i_025    tia_h_in_001_015-    120831.44397548852
Rh001_026_015+    i_026    tia_h_in_001_015+    5000
Rh001_026_015-    i_026    tia_h_in_001_015-    80511.3256230622
Rh001_027_015+    i_027    tia_h_in_001_015+    120864.63601072058
Rh001_027_015-    i_027    tia_h_in_001_015-    80795.6451005659
Rh001_028_015+    i_028    tia_h_in_001_015+    72851.58940478401
Rh001_028_015-    i_028    tia_h_in_001_015-    119302.97667044237
Rh001_029_015+    i_029    tia_h_in_001_015+    122141.30073896536
Rh001_029_015-    i_029    tia_h_in_001_015-    76661.14179843181
Rh001_030_015+    i_030    tia_h_in_001_015+    119271.47333271494
Rh001_030_015-    i_030    tia_h_in_001_015-    97021.04199301725
Rh001_031_015+    i_031    tia_h_in_001_015+    58104.96024857979
Rh001_031_015-    i_031    tia_h_in_001_015-    119902.98355165585
Rh001_032_015+    i_032    tia_h_in_001_015+    118075.50096856373
Rh001_032_015-    i_032    tia_h_in_001_015-    75280.13978785997
Rh001_033_015+    i_033    tia_h_in_001_015+    120584.47981618161
Rh001_033_015-    i_033    tia_h_in_001_015-    60955.68290138255
Rh001_034_015+    i_034    tia_h_in_001_015+    120636.48116671642
Rh001_034_015-    i_034    tia_h_in_001_015-    66386.50285627852
Rh001_035_015+    i_035    tia_h_in_001_015+    120087.44256993911
Rh001_035_015-    i_035    tia_h_in_001_015-    84137.11596610055
Rh001_036_015+    i_036    tia_h_in_001_015+    119805.85514208721
Rh001_036_015-    i_036    tia_h_in_001_015-    70627.55233864371
Rh001_037_015+    i_037    tia_h_in_001_015+    121276.95374337304
Rh001_037_015-    i_037    tia_h_in_001_015-    5000
Rh001_038_015+    i_038    tia_h_in_001_015+    85870.224988958
Rh001_038_015-    i_038    tia_h_in_001_015-    120332.19931302119
Rh001_039_015+    i_039    tia_h_in_001_015+    107587.15254050354
Rh001_039_015-    i_039    tia_h_in_001_015-    120120.37302899513
Rh001_040_015+    i_040    tia_h_in_001_015+    120192.55778710131
Rh001_040_015-    i_040    tia_h_in_001_015-    79733.46005192983
Rh001_041_015+    i_041    tia_h_in_001_015+    121607.73501361054
Rh001_041_015-    i_041    tia_h_in_001_015-    59058.03507034096
Rh001_042_015+    i_042    tia_h_in_001_015+    120512.46816093232
Rh001_042_015-    i_042    tia_h_in_001_015-    79719.65640027977
Rh001_043_015+    i_043    tia_h_in_001_015+    120171.99415897732
Rh001_043_015-    i_043    tia_h_in_001_015-    74484.9970605876
Rh001_044_015+    i_044    tia_h_in_001_015+    119511.91374399603
Rh001_044_015-    i_044    tia_h_in_001_015-    80073.61420572147
Rh001_045_015+    i_045    tia_h_in_001_015+    119380.58678161324
Rh001_045_015-    i_045    tia_h_in_001_015-    54283.83309567027
Rh001_046_015+    i_046    tia_h_in_001_015+    104834.53111067195
Rh001_046_015-    i_046    tia_h_in_001_015-    118983.73356872889
Rh001_047_015+    i_047    tia_h_in_001_015+    119907.97097466607
Rh001_047_015-    i_047    tia_h_in_001_015-    60454.66449663913
Rh001_048_015+    i_048    tia_h_in_001_015+    120000
Rh001_048_015-    i_048    tia_h_in_001_015-    57209.04761200684
Rh001_049_015+    i_049    tia_h_in_001_015+    121067.8997152489
Rh001_049_015-    i_049    tia_h_in_001_015-    56885.214751399806
Rh001_050_015+    i_050    tia_h_in_001_015+    120000
Rh001_050_015-    i_050    tia_h_in_001_015-    120462.10160297914
Rh001_051_015+    i_051    tia_h_in_001_015+    118807.20292121699
Rh001_051_015-    i_051    tia_h_in_001_015-    65544.89300762562
Rh001_052_015+    i_052    tia_h_in_001_015+    121654.28294041626
Rh001_052_015-    i_052    tia_h_in_001_015-    74327.16293795544
Rh001_053_015+    i_053    tia_h_in_001_015+    63733.287858010524
Rh001_053_015-    i_053    tia_h_in_001_015-    121720.09756678491
Rh001_054_015+    i_054    tia_h_in_001_015+    77911.60418448251
Rh001_054_015-    i_054    tia_h_in_001_015-    117642.8636320814
Rh001_055_015+    i_055    tia_h_in_001_015+    74541.69794204795
Rh001_055_015-    i_055    tia_h_in_001_015-    120933.71860280272
Rh001_056_015+    i_056    tia_h_in_001_015+    120826.87714095219
Rh001_056_015-    i_056    tia_h_in_001_015-    52756.99839794678
Rh001_057_015+    i_057    tia_h_in_001_015+    5000
Rh001_057_015-    i_057    tia_h_in_001_015-    5000
Rh001_058_015+    i_058    tia_h_in_001_015+    118919.51938352906
Rh001_058_015-    i_058    tia_h_in_001_015-    75934.38969855173
Rh001_059_015+    i_059    tia_h_in_001_015+    62804.48641094691
Rh001_059_015-    i_059    tia_h_in_001_015-    120497.02882180734
Rh001_060_015+    i_060    tia_h_in_001_015+    113984.38449101105
Rh001_060_015-    i_060    tia_h_in_001_015-    118095.93010197341
Rh001_061_015+    i_061    tia_h_in_001_015+    117965.23814118399
Rh001_061_015-    i_061    tia_h_in_001_015-    59669.77662109178
Rh001_062_015+    i_062    tia_h_in_001_015+    5000
Rh001_062_015-    i_062    tia_h_in_001_015-    106682.62461399045
Rh001_063_015+    i_063    tia_h_in_001_015+    120000
Rh001_063_015-    i_063    tia_h_in_001_015-    56780.10863072095
Rh001_064_015+    i_064    tia_h_in_001_015+    120720.6721752781
Rh001_064_015-    i_064    tia_h_in_001_015-    90665.72413302884

* Neuron 16
Rh001_001_016+    i_001    tia_h_in_001_016+    27832.532207571097
Rh001_001_016-    i_001    tia_h_in_001_016-    119697.45766816757
Rh001_002_016+    i_002    tia_h_in_001_016+    25139.673620763817
Rh001_002_016-    i_002    tia_h_in_001_016-    120000
Rh001_003_016+    i_003    tia_h_in_001_016+    77730.51232181903
Rh001_003_016-    i_003    tia_h_in_001_016-    120815.23234705371
Rh001_004_016+    i_004    tia_h_in_001_016+    120000
Rh001_004_016-    i_004    tia_h_in_001_016-    42878.3187586264
Rh001_005_016+    i_005    tia_h_in_001_016+    120524.30936946908
Rh001_005_016-    i_005    tia_h_in_001_016-    20519.215487499278
Rh001_006_016+    i_006    tia_h_in_001_016+    120410.26662432449
Rh001_006_016-    i_006    tia_h_in_001_016-    17901.800620648202
Rh001_007_016+    i_007    tia_h_in_001_016+    119791.4229761061
Rh001_007_016-    i_007    tia_h_in_001_016-    95759.93080919914
Rh001_008_016+    i_008    tia_h_in_001_016+    5000
Rh001_008_016-    i_008    tia_h_in_001_016-    120565.93052510085
Rh001_009_016+    i_009    tia_h_in_001_016+    120358.21600979
Rh001_009_016-    i_009    tia_h_in_001_016-    66633.5665945886
Rh001_010_016+    i_010    tia_h_in_001_016+    119554.81044770498
Rh001_010_016-    i_010    tia_h_in_001_016-    120000
Rh001_011_016+    i_011    tia_h_in_001_016+    121093.71712761588
Rh001_011_016-    i_011    tia_h_in_001_016-    48068.98210689664
Rh001_012_016+    i_012    tia_h_in_001_016+    120425.71360471561
Rh001_012_016-    i_012    tia_h_in_001_016-    44647.14709507756
Rh001_013_016+    i_013    tia_h_in_001_016+    119538.62746559293
Rh001_013_016-    i_013    tia_h_in_001_016-    84072.68517401641
Rh001_014_016+    i_014    tia_h_in_001_016+    89156.21854419008
Rh001_014_016-    i_014    tia_h_in_001_016-    120651.66764214588
Rh001_015_016+    i_015    tia_h_in_001_016+    120000
Rh001_015_016-    i_015    tia_h_in_001_016-    120337.25725928388
Rh001_016_016+    i_016    tia_h_in_001_016+    39809.87585951941
Rh001_016_016-    i_016    tia_h_in_001_016-    121169.19371909916
Rh001_017_016+    i_017    tia_h_in_001_016+    121554.25279198555
Rh001_017_016-    i_017    tia_h_in_001_016-    104676.59069506623
Rh001_018_016+    i_018    tia_h_in_001_016+    44379.326543846066
Rh001_018_016-    i_018    tia_h_in_001_016-    120000
Rh001_019_016+    i_019    tia_h_in_001_016+    119649.23471543979
Rh001_019_016-    i_019    tia_h_in_001_016-    97668.17244827143
Rh001_020_016+    i_020    tia_h_in_001_016+    5000
Rh001_020_016-    i_020    tia_h_in_001_016-    49165.38879378579
Rh001_021_016+    i_021    tia_h_in_001_016+    120442.76576516968
Rh001_021_016-    i_021    tia_h_in_001_016-    34420.62002803935
Rh001_022_016+    i_022    tia_h_in_001_016+    121387.07088968105
Rh001_022_016-    i_022    tia_h_in_001_016-    116703.20212010869
Rh001_023_016+    i_023    tia_h_in_001_016+    120861.98543885656
Rh001_023_016-    i_023    tia_h_in_001_016-    61172.22430171714
Rh001_024_016+    i_024    tia_h_in_001_016+    5000
Rh001_024_016-    i_024    tia_h_in_001_016-    120494.77038652434
Rh001_025_016+    i_025    tia_h_in_001_016+    5000
Rh001_025_016-    i_025    tia_h_in_001_016-    120659.62014179178
Rh001_026_016+    i_026    tia_h_in_001_016+    119535.0126253259
Rh001_026_016-    i_026    tia_h_in_001_016-    62405.84048547506
Rh001_027_016+    i_027    tia_h_in_001_016+    121383.51661924145
Rh001_027_016-    i_027    tia_h_in_001_016-    66454.85954657022
Rh001_028_016+    i_028    tia_h_in_001_016+    119451.04199662602
Rh001_028_016-    i_028    tia_h_in_001_016-    89264.59147148787
Rh001_029_016+    i_029    tia_h_in_001_016+    117327.29340663138
Rh001_029_016-    i_029    tia_h_in_001_016-    120256.09227688774
Rh001_030_016+    i_030    tia_h_in_001_016+    119508.21348361508
Rh001_030_016-    i_030    tia_h_in_001_016-    89329.25660533253
Rh001_031_016+    i_031    tia_h_in_001_016+    48830.11105452216
Rh001_031_016-    i_031    tia_h_in_001_016-    120770.30060795548
Rh001_032_016+    i_032    tia_h_in_001_016+    57254.401389684535
Rh001_032_016-    i_032    tia_h_in_001_016-    120571.84752511942
Rh001_033_016+    i_033    tia_h_in_001_016+    116089.58632857156
Rh001_033_016-    i_033    tia_h_in_001_016-    118537.10805470741
Rh001_034_016+    i_034    tia_h_in_001_016+    112084.13551933097
Rh001_034_016-    i_034    tia_h_in_001_016-    119060.47304633704
Rh001_035_016+    i_035    tia_h_in_001_016+    119760.96810701405
Rh001_035_016-    i_035    tia_h_in_001_016-    43821.666990002224
Rh001_036_016+    i_036    tia_h_in_001_016+    119337.57451032902
Rh001_036_016-    i_036    tia_h_in_001_016-    37912.54703089404
Rh001_037_016+    i_037    tia_h_in_001_016+    74940.04530965016
Rh001_037_016-    i_037    tia_h_in_001_016-    119588.11696283211
Rh001_038_016+    i_038    tia_h_in_001_016+    36784.90905931099
Rh001_038_016-    i_038    tia_h_in_001_016-    119721.05485503355
Rh001_039_016+    i_039    tia_h_in_001_016+    79548.90757777216
Rh001_039_016-    i_039    tia_h_in_001_016-    120202.08740972544
Rh001_040_016+    i_040    tia_h_in_001_016+    41291.89121711025
Rh001_040_016-    i_040    tia_h_in_001_016-    120091.82419991055
Rh001_041_016+    i_041    tia_h_in_001_016+    120858.30760426327
Rh001_041_016-    i_041    tia_h_in_001_016-    44328.95132061535
Rh001_042_016+    i_042    tia_h_in_001_016+    119977.45282153478
Rh001_042_016-    i_042    tia_h_in_001_016-    60987.431806998175
Rh001_043_016+    i_043    tia_h_in_001_016+    119773.96833089308
Rh001_043_016-    i_043    tia_h_in_001_016-    5000
Rh001_044_016+    i_044    tia_h_in_001_016+    39735.50872290538
Rh001_044_016-    i_044    tia_h_in_001_016-    118779.28668828002
Rh001_045_016+    i_045    tia_h_in_001_016+    37242.92331430243
Rh001_045_016-    i_045    tia_h_in_001_016-    121128.19235051771
Rh001_046_016+    i_046    tia_h_in_001_016+    43005.08876592589
Rh001_046_016-    i_046    tia_h_in_001_016-    118823.07473266071
Rh001_047_016+    i_047    tia_h_in_001_016+    70668.20390884536
Rh001_047_016-    i_047    tia_h_in_001_016-    118547.57889439503
Rh001_048_016+    i_048    tia_h_in_001_016+    118774.13790415674
Rh001_048_016-    i_048    tia_h_in_001_016-    39983.732844926555
Rh001_049_016+    i_049    tia_h_in_001_016+    120000
Rh001_049_016-    i_049    tia_h_in_001_016-    5000
Rh001_050_016+    i_050    tia_h_in_001_016+    119844.22293617755
Rh001_050_016-    i_050    tia_h_in_001_016-    40837.68217746429
Rh001_051_016+    i_051    tia_h_in_001_016+    121504.07338487516
Rh001_051_016-    i_051    tia_h_in_001_016-    50417.942417929415
Rh001_052_016+    i_052    tia_h_in_001_016+    56681.6146912795
Rh001_052_016-    i_052    tia_h_in_001_016-    119613.21197825935
Rh001_053_016+    i_053    tia_h_in_001_016+    51473.65902540904
Rh001_053_016-    i_053    tia_h_in_001_016-    120193.53104244267
Rh001_054_016+    i_054    tia_h_in_001_016+    31238.9762698155
Rh001_054_016-    i_054    tia_h_in_001_016-    118718.3170404038
Rh001_055_016+    i_055    tia_h_in_001_016+    52766.089426330065
Rh001_055_016-    i_055    tia_h_in_001_016-    120000
Rh001_056_016+    i_056    tia_h_in_001_016+    120257.17095610207
Rh001_056_016-    i_056    tia_h_in_001_016-    57615.156001581694
Rh001_057_016+    i_057    tia_h_in_001_016+    121258.02021157918
Rh001_057_016-    i_057    tia_h_in_001_016-    41533.07249035249
Rh001_058_016+    i_058    tia_h_in_001_016+    119604.48347012646
Rh001_058_016-    i_058    tia_h_in_001_016-    63628.38846567681
Rh001_059_016+    i_059    tia_h_in_001_016+    27774.592526255215
Rh001_059_016-    i_059    tia_h_in_001_016-    120000
Rh001_060_016+    i_060    tia_h_in_001_016+    22919.06954564759
Rh001_060_016-    i_060    tia_h_in_001_016-    119736.69890960421
Rh001_061_016+    i_061    tia_h_in_001_016+    25164.876502334155
Rh001_061_016-    i_061    tia_h_in_001_016-    120769.37366023328
Rh001_062_016+    i_062    tia_h_in_001_016+    120525.63329511815
Rh001_062_016-    i_062    tia_h_in_001_016-    99501.85140368382
Rh001_063_016+    i_063    tia_h_in_001_016+    120225.93420869844
Rh001_063_016-    i_063    tia_h_in_001_016-    25735.14290021918
Rh001_064_016+    i_064    tia_h_in_001_016+    120000
Rh001_064_016-    i_064    tia_h_in_001_016-    24509.674874361757

* Neuron 17
Rh001_001_017+    i_001    tia_h_in_001_017+    118794.93472202236
Rh001_001_017-    i_001    tia_h_in_001_017-    46827.03837072743
Rh001_002_017+    i_002    tia_h_in_001_017+    77616.85456879552
Rh001_002_017-    i_002    tia_h_in_001_017-    119354.16130196121
Rh001_003_017+    i_003    tia_h_in_001_017+    120267.25844598767
Rh001_003_017-    i_003    tia_h_in_001_017-    30536.080085438258
Rh001_004_017+    i_004    tia_h_in_001_017+    119654.94247541875
Rh001_004_017-    i_004    tia_h_in_001_017-    13641.621089824286
Rh001_005_017+    i_005    tia_h_in_001_017+    120342.31815112715
Rh001_005_017-    i_005    tia_h_in_001_017-    120000
Rh001_006_017+    i_006    tia_h_in_001_017+    36972.70142529555
Rh001_006_017-    i_006    tia_h_in_001_017-    120093.81438670009
Rh001_007_017+    i_007    tia_h_in_001_017+    31129.43113874689
Rh001_007_017-    i_007    tia_h_in_001_017-    120000
Rh001_008_017+    i_008    tia_h_in_001_017+    31464.360413496783
Rh001_008_017-    i_008    tia_h_in_001_017-    120391.48982539053
Rh001_009_017+    i_009    tia_h_in_001_017+    121267.92175518256
Rh001_009_017-    i_009    tia_h_in_001_017-    71814.34656831341
Rh001_010_017+    i_010    tia_h_in_001_017+    118311.3280671651
Rh001_010_017-    i_010    tia_h_in_001_017-    41586.57145263021
Rh001_011_017+    i_011    tia_h_in_001_017+    119886.12055644112
Rh001_011_017-    i_011    tia_h_in_001_017-    5000
Rh001_012_017+    i_012    tia_h_in_001_017+    118604.43157528946
Rh001_012_017-    i_012    tia_h_in_001_017-    51457.6517738974
Rh001_013_017+    i_013    tia_h_in_001_017+    53836.28716834618
Rh001_013_017-    i_013    tia_h_in_001_017-    120571.13139083944
Rh001_014_017+    i_014    tia_h_in_001_017+    23725.75131916746
Rh001_014_017-    i_014    tia_h_in_001_017-    119662.08843036005
Rh001_015_017+    i_015    tia_h_in_001_017+    75372.10603041032
Rh001_015_017-    i_015    tia_h_in_001_017-    118856.39760029534
Rh001_016_017+    i_016    tia_h_in_001_017+    119280.19658695953
Rh001_016_017-    i_016    tia_h_in_001_017-    94378.55878734187
Rh001_017_017+    i_017    tia_h_in_001_017+    119171.89280360797
Rh001_017_017-    i_017    tia_h_in_001_017-    81797.22011740366
Rh001_018_017+    i_018    tia_h_in_001_017+    119435.3716571852
Rh001_018_017-    i_018    tia_h_in_001_017-    5000
Rh001_019_017+    i_019    tia_h_in_001_017+    121187.23385977732
Rh001_019_017-    i_019    tia_h_in_001_017-    33774.02837559075
Rh001_020_017+    i_020    tia_h_in_001_017+    120631.50491859566
Rh001_020_017-    i_020    tia_h_in_001_017-    100616.36914558308
Rh001_021_017+    i_021    tia_h_in_001_017+    43613.17661542547
Rh001_021_017-    i_021    tia_h_in_001_017-    120438.23305199621
Rh001_022_017+    i_022    tia_h_in_001_017+    62620.597872909544
Rh001_022_017-    i_022    tia_h_in_001_017-    118991.10565528338
Rh001_023_017+    i_023    tia_h_in_001_017+    51008.00410661321
Rh001_023_017-    i_023    tia_h_in_001_017-    121791.99221966266
Rh001_024_017+    i_024    tia_h_in_001_017+    119184.59474262585
Rh001_024_017-    i_024    tia_h_in_001_017-    49332.554388167075
Rh001_025_017+    i_025    tia_h_in_001_017+    78268.13581260518
Rh001_025_017-    i_025    tia_h_in_001_017-    120000
Rh001_026_017+    i_026    tia_h_in_001_017+    78285.02541391207
Rh001_026_017-    i_026    tia_h_in_001_017-    119487.12974831539
Rh001_027_017+    i_027    tia_h_in_001_017+    53029.43705093152
Rh001_027_017-    i_027    tia_h_in_001_017-    121149.90581291256
Rh001_028_017+    i_028    tia_h_in_001_017+    31225.99398199212
Rh001_028_017-    i_028    tia_h_in_001_017-    119817.12222909502
Rh001_029_017+    i_029    tia_h_in_001_017+    19438.06609107247
Rh001_029_017-    i_029    tia_h_in_001_017-    121104.79393465983
Rh001_030_017+    i_030    tia_h_in_001_017+    38937.61488905819
Rh001_030_017-    i_030    tia_h_in_001_017-    120821.35135550665
Rh001_031_017+    i_031    tia_h_in_001_017+    120377.25073316443
Rh001_031_017-    i_031    tia_h_in_001_017-    30500.837805292475
Rh001_032_017+    i_032    tia_h_in_001_017+    120588.12835747434
Rh001_032_017-    i_032    tia_h_in_001_017-    62590.04891230923
Rh001_033_017+    i_033    tia_h_in_001_017+    119293.54445871226
Rh001_033_017-    i_033    tia_h_in_001_017-    74091.69274106219
Rh001_034_017+    i_034    tia_h_in_001_017+    118530.46072833185
Rh001_034_017-    i_034    tia_h_in_001_017-    27349.634365782236
Rh001_035_017+    i_035    tia_h_in_001_017+    27633.64717223433
Rh001_035_017-    i_035    tia_h_in_001_017-    119923.32848335218
Rh001_036_017+    i_036    tia_h_in_001_017+    21719.976515520946
Rh001_036_017-    i_036    tia_h_in_001_017-    121687.43059166783
Rh001_037_017+    i_037    tia_h_in_001_017+    5000
Rh001_037_017-    i_037    tia_h_in_001_017-    120191.64701528076
Rh001_038_017+    i_038    tia_h_in_001_017+    71968.29009058615
Rh001_038_017-    i_038    tia_h_in_001_017-    119606.26173516139
Rh001_039_017+    i_039    tia_h_in_001_017+    119991.35790456632
Rh001_039_017-    i_039    tia_h_in_001_017-    73158.4472374898
Rh001_040_017+    i_040    tia_h_in_001_017+    57338.87132166247
Rh001_040_017-    i_040    tia_h_in_001_017-    120000
Rh001_041_017+    i_041    tia_h_in_001_017+    69671.26024170626
Rh001_041_017-    i_041    tia_h_in_001_017-    120136.53705615514
Rh001_042_017+    i_042    tia_h_in_001_017+    49546.66471749548
Rh001_042_017-    i_042    tia_h_in_001_017-    119652.32781501966
Rh001_043_017+    i_043    tia_h_in_001_017+    5000
Rh001_043_017-    i_043    tia_h_in_001_017-    118472.91783440998
Rh001_044_017+    i_044    tia_h_in_001_017+    70089.10440819604
Rh001_044_017-    i_044    tia_h_in_001_017-    120000
Rh001_045_017+    i_045    tia_h_in_001_017+    120526.46310980644
Rh001_045_017-    i_045    tia_h_in_001_017-    120000
Rh001_046_017+    i_046    tia_h_in_001_017+    119431.94613246771
Rh001_046_017-    i_046    tia_h_in_001_017-    120000
Rh001_047_017+    i_047    tia_h_in_001_017+    117906.11220862839
Rh001_047_017-    i_047    tia_h_in_001_017-    68313.86195044016
Rh001_048_017+    i_048    tia_h_in_001_017+    120266.60655490063
Rh001_048_017-    i_048    tia_h_in_001_017-    107308.84398205052
Rh001_049_017+    i_049    tia_h_in_001_017+    119380.10239089593
Rh001_049_017-    i_049    tia_h_in_001_017-    56158.94050902814
Rh001_050_017+    i_050    tia_h_in_001_017+    5000
Rh001_050_017-    i_050    tia_h_in_001_017-    119139.61945224911
Rh001_051_017+    i_051    tia_h_in_001_017+    41313.74002435476
Rh001_051_017-    i_051    tia_h_in_001_017-    120000
Rh001_052_017+    i_052    tia_h_in_001_017+    45344.1518131135
Rh001_052_017-    i_052    tia_h_in_001_017-    118716.77077752782
Rh001_053_017+    i_053    tia_h_in_001_017+    119370.95780216841
Rh001_053_017-    i_053    tia_h_in_001_017-    68446.40815212505
Rh001_054_017+    i_054    tia_h_in_001_017+    120068.78578159971
Rh001_054_017-    i_054    tia_h_in_001_017-    26396.512630377074
Rh001_055_017+    i_055    tia_h_in_001_017+    120720.83924134493
Rh001_055_017-    i_055    tia_h_in_001_017-    51898.76037310404
Rh001_056_017+    i_056    tia_h_in_001_017+    120653.63791483454
Rh001_056_017-    i_056    tia_h_in_001_017-    39278.228090785655
Rh001_057_017+    i_057    tia_h_in_001_017+    41770.55471712812
Rh001_057_017-    i_057    tia_h_in_001_017-    118368.2043936838
Rh001_058_017+    i_058    tia_h_in_001_017+    32184.592059415747
Rh001_058_017-    i_058    tia_h_in_001_017-    119417.19019282375
Rh001_059_017+    i_059    tia_h_in_001_017+    35727.58138190437
Rh001_059_017-    i_059    tia_h_in_001_017-    5000
Rh001_060_017+    i_060    tia_h_in_001_017+    121863.12461706983
Rh001_060_017-    i_060    tia_h_in_001_017-    32219.926067620407
Rh001_061_017+    i_061    tia_h_in_001_017+    118497.9215835261
Rh001_061_017-    i_061    tia_h_in_001_017-    14451.354369328386
Rh001_062_017+    i_062    tia_h_in_001_017+    120392.65661609638
Rh001_062_017-    i_062    tia_h_in_001_017-    32604.582954338162
Rh001_063_017+    i_063    tia_h_in_001_017+    57419.41277049883
Rh001_063_017-    i_063    tia_h_in_001_017-    119560.5200191886
Rh001_064_017+    i_064    tia_h_in_001_017+    101587.53808096051
Rh001_064_017-    i_064    tia_h_in_001_017-    119534.66123163869

* Neuron 18
Rh001_001_018+    i_001    tia_h_in_001_018+    119266.59229089631
Rh001_001_018-    i_001    tia_h_in_001_018-    30698.993641953133
Rh001_002_018+    i_002    tia_h_in_001_018+    120563.18939454012
Rh001_002_018-    i_002    tia_h_in_001_018-    28785.436012641825
Rh001_003_018+    i_003    tia_h_in_001_018+    119611.33955950796
Rh001_003_018-    i_003    tia_h_in_001_018-    75446.31184313587
Rh001_004_018+    i_004    tia_h_in_001_018+    119332.01616492696
Rh001_004_018-    i_004    tia_h_in_001_018-    120000
Rh001_005_018+    i_005    tia_h_in_001_018+    115721.93108456547
Rh001_005_018-    i_005    tia_h_in_001_018-    121673.78145109503
Rh001_006_018+    i_006    tia_h_in_001_018+    120453.7802629931
Rh001_006_018-    i_006    tia_h_in_001_018-    62292.99415432728
Rh001_007_018+    i_007    tia_h_in_001_018+    82922.95469174683
Rh001_007_018-    i_007    tia_h_in_001_018-    120083.37626638582
Rh001_008_018+    i_008    tia_h_in_001_018+    55643.007595975236
Rh001_008_018-    i_008    tia_h_in_001_018-    120000
Rh001_009_018+    i_009    tia_h_in_001_018+    120478.70370654354
Rh001_009_018-    i_009    tia_h_in_001_018-    36952.67519871133
Rh001_010_018+    i_010    tia_h_in_001_018+    119834.0804819477
Rh001_010_018-    i_010    tia_h_in_001_018-    5000
Rh001_011_018+    i_011    tia_h_in_001_018+    61489.045387247184
Rh001_011_018-    i_011    tia_h_in_001_018-    120000
Rh001_012_018+    i_012    tia_h_in_001_018+    61626.488851848204
Rh001_012_018-    i_012    tia_h_in_001_018-    120420.16041965547
Rh001_013_018+    i_013    tia_h_in_001_018+    5000
Rh001_013_018-    i_013    tia_h_in_001_018-    107057.77483747306
Rh001_014_018+    i_014    tia_h_in_001_018+    57415.18420265447
Rh001_014_018-    i_014    tia_h_in_001_018-    119114.5511431548
Rh001_015_018+    i_015    tia_h_in_001_018+    67996.46020939096
Rh001_015_018-    i_015    tia_h_in_001_018-    119533.44065608774
Rh001_016_018+    i_016    tia_h_in_001_018+    117584.00795394398
Rh001_016_018-    i_016    tia_h_in_001_018-    47745.70608624806
Rh001_017_018+    i_017    tia_h_in_001_018+    89671.35269154742
Rh001_017_018-    i_017    tia_h_in_001_018-    118281.45150046704
Rh001_018_018+    i_018    tia_h_in_001_018+    72899.22646574961
Rh001_018_018-    i_018    tia_h_in_001_018-    120341.93464077915
Rh001_019_018+    i_019    tia_h_in_001_018+    5000
Rh001_019_018-    i_019    tia_h_in_001_018-    120783.60805679884
Rh001_020_018+    i_020    tia_h_in_001_018+    121526.12347811522
Rh001_020_018-    i_020    tia_h_in_001_018-    62723.83772832352
Rh001_021_018+    i_021    tia_h_in_001_018+    79303.25540639537
Rh001_021_018-    i_021    tia_h_in_001_018-    122415.72343864117
Rh001_022_018+    i_022    tia_h_in_001_018+    120118.69451468816
Rh001_022_018-    i_022    tia_h_in_001_018-    106411.53070683783
Rh001_023_018+    i_023    tia_h_in_001_018+    118627.45993930985
Rh001_023_018-    i_023    tia_h_in_001_018-    85653.90876766539
Rh001_024_018+    i_024    tia_h_in_001_018+    102697.04592064144
Rh001_024_018-    i_024    tia_h_in_001_018-    117906.63786004063
Rh001_025_018+    i_025    tia_h_in_001_018+    64940.29926143623
Rh001_025_018-    i_025    tia_h_in_001_018-    119455.4404910485
Rh001_026_018+    i_026    tia_h_in_001_018+    44449.88279520814
Rh001_026_018-    i_026    tia_h_in_001_018-    119720.99176983704
Rh001_027_018+    i_027    tia_h_in_001_018+    5000
Rh001_027_018-    i_027    tia_h_in_001_018-    119781.15826998027
Rh001_028_018+    i_028    tia_h_in_001_018+    53849.72802171319
Rh001_028_018-    i_028    tia_h_in_001_018-    120200.66645285695
Rh001_029_018+    i_029    tia_h_in_001_018+    119763.24985709516
Rh001_029_018-    i_029    tia_h_in_001_018-    48700.242791054254
Rh001_030_018+    i_030    tia_h_in_001_018+    120177.03717484807
Rh001_030_018-    i_030    tia_h_in_001_018-    44919.56890488154
Rh001_031_018+    i_031    tia_h_in_001_018+    44826.72776671601
Rh001_031_018-    i_031    tia_h_in_001_018-    119659.55499033391
Rh001_032_018+    i_032    tia_h_in_001_018+    119718.16007611617
Rh001_032_018-    i_032    tia_h_in_001_018-    95358.55243372497
Rh001_033_018+    i_033    tia_h_in_001_018+    35184.00813725485
Rh001_033_018-    i_033    tia_h_in_001_018-    118957.92262123681
Rh001_034_018+    i_034    tia_h_in_001_018+    53765.567900034046
Rh001_034_018-    i_034    tia_h_in_001_018-    120990.89626922672
Rh001_035_018+    i_035    tia_h_in_001_018+    119614.51775923611
Rh001_035_018-    i_035    tia_h_in_001_018-    81490.66936282332
Rh001_036_018+    i_036    tia_h_in_001_018+    65901.13339539045
Rh001_036_018-    i_036    tia_h_in_001_018-    121029.81905798506
Rh001_037_018+    i_037    tia_h_in_001_018+    120000
Rh001_037_018-    i_037    tia_h_in_001_018-    120804.7936667826
Rh001_038_018+    i_038    tia_h_in_001_018+    47918.115041238256
Rh001_038_018-    i_038    tia_h_in_001_018-    120000
Rh001_039_018+    i_039    tia_h_in_001_018+    63099.69035965014
Rh001_039_018-    i_039    tia_h_in_001_018-    120651.11494161005
Rh001_040_018+    i_040    tia_h_in_001_018+    22850.837613978652
Rh001_040_018-    i_040    tia_h_in_001_018-    118586.16410816864
Rh001_041_018+    i_041    tia_h_in_001_018+    119379.0495191284
Rh001_041_018-    i_041    tia_h_in_001_018-    78653.40681512794
Rh001_042_018+    i_042    tia_h_in_001_018+    119649.4724555453
Rh001_042_018-    i_042    tia_h_in_001_018-    62802.39595973425
Rh001_043_018+    i_043    tia_h_in_001_018+    119544.15088120039
Rh001_043_018-    i_043    tia_h_in_001_018-    101450.45191486014
Rh001_044_018+    i_044    tia_h_in_001_018+    118334.37785970363
Rh001_044_018-    i_044    tia_h_in_001_018-    118876.00376825673
Rh001_045_018+    i_045    tia_h_in_001_018+    119139.16206874234
Rh001_045_018-    i_045    tia_h_in_001_018-    84777.4928590408
Rh001_046_018+    i_046    tia_h_in_001_018+    34298.239488398845
Rh001_046_018-    i_046    tia_h_in_001_018-    5000
Rh001_047_018+    i_047    tia_h_in_001_018+    45672.40604154794
Rh001_047_018-    i_047    tia_h_in_001_018-    120244.70036410102
Rh001_048_018+    i_048    tia_h_in_001_018+    35720.145294525726
Rh001_048_018-    i_048    tia_h_in_001_018-    119623.37898268056
Rh001_049_018+    i_049    tia_h_in_001_018+    118395.86209180945
Rh001_049_018-    i_049    tia_h_in_001_018-    92089.12992840893
Rh001_050_018+    i_050    tia_h_in_001_018+    98993.13043796479
Rh001_050_018-    i_050    tia_h_in_001_018-    120941.11172949994
Rh001_051_018+    i_051    tia_h_in_001_018+    119420.033216115
Rh001_051_018-    i_051    tia_h_in_001_018-    79286.69691939598
Rh001_052_018+    i_052    tia_h_in_001_018+    120216.69080243903
Rh001_052_018-    i_052    tia_h_in_001_018-    70957.57180113916
Rh001_053_018+    i_053    tia_h_in_001_018+    120560.1758301777
Rh001_053_018-    i_053    tia_h_in_001_018-    90122.96127674544
Rh001_054_018+    i_054    tia_h_in_001_018+    118610.07005356568
Rh001_054_018-    i_054    tia_h_in_001_018-    63719.6492335011
Rh001_055_018+    i_055    tia_h_in_001_018+    71143.08326931314
Rh001_055_018-    i_055    tia_h_in_001_018-    118662.42181873461
Rh001_056_018+    i_056    tia_h_in_001_018+    121614.69827339864
Rh001_056_018-    i_056    tia_h_in_001_018-    21678.186290900987
Rh001_057_018+    i_057    tia_h_in_001_018+    67616.19752190566
Rh001_057_018-    i_057    tia_h_in_001_018-    5000
Rh001_058_018+    i_058    tia_h_in_001_018+    93940.28223038075
Rh001_058_018-    i_058    tia_h_in_001_018-    121399.11335845539
Rh001_059_018+    i_059    tia_h_in_001_018+    119036.3299027612
Rh001_059_018-    i_059    tia_h_in_001_018-    73691.56331997836
Rh001_060_018+    i_060    tia_h_in_001_018+    44403.82522450149
Rh001_060_018-    i_060    tia_h_in_001_018-    118366.19750634962
Rh001_061_018+    i_061    tia_h_in_001_018+    120746.15444896273
Rh001_061_018-    i_061    tia_h_in_001_018-    74406.27128927871
Rh001_062_018+    i_062    tia_h_in_001_018+    120653.09938059845
Rh001_062_018-    i_062    tia_h_in_001_018-    47736.81307485108
Rh001_063_018+    i_063    tia_h_in_001_018+    121293.86731299976
Rh001_063_018-    i_063    tia_h_in_001_018-    17273.29016772587
Rh001_064_018+    i_064    tia_h_in_001_018+    5000
Rh001_064_018-    i_064    tia_h_in_001_018-    24481.400916449635

* Neuron 19
Rh001_001_019+    i_001    tia_h_in_001_019+    120000
Rh001_001_019-    i_001    tia_h_in_001_019-    120831.76223418185
Rh001_002_019+    i_002    tia_h_in_001_019+    48866.470780955264
Rh001_002_019-    i_002    tia_h_in_001_019-    119482.57353271067
Rh001_003_019+    i_003    tia_h_in_001_019+    20859.9765444617
Rh001_003_019-    i_003    tia_h_in_001_019-    120603.72023724423
Rh001_004_019+    i_004    tia_h_in_001_019+    79244.48736126848
Rh001_004_019-    i_004    tia_h_in_001_019-    121184.38479067099
Rh001_005_019+    i_005    tia_h_in_001_019+    121036.15814809313
Rh001_005_019-    i_005    tia_h_in_001_019-    39877.09936014656
Rh001_006_019+    i_006    tia_h_in_001_019+    120000
Rh001_006_019-    i_006    tia_h_in_001_019-    29981.035294472378
Rh001_007_019+    i_007    tia_h_in_001_019+    120000
Rh001_007_019-    i_007    tia_h_in_001_019-    120000
Rh001_008_019+    i_008    tia_h_in_001_019+    118384.66036477016
Rh001_008_019-    i_008    tia_h_in_001_019-    39825.85207128536
Rh001_009_019+    i_009    tia_h_in_001_019+    70254.81752550919
Rh001_009_019-    i_009    tia_h_in_001_019-    120207.2160398045
Rh001_010_019+    i_010    tia_h_in_001_019+    38337.137671052005
Rh001_010_019-    i_010    tia_h_in_001_019-    120012.44472189325
Rh001_011_019+    i_011    tia_h_in_001_019+    119403.9048916423
Rh001_011_019-    i_011    tia_h_in_001_019-    70431.71174253825
Rh001_012_019+    i_012    tia_h_in_001_019+    119611.58939170564
Rh001_012_019-    i_012    tia_h_in_001_019-    5000
Rh001_013_019+    i_013    tia_h_in_001_019+    119778.79036103033
Rh001_013_019-    i_013    tia_h_in_001_019-    46859.638101624885
Rh001_014_019+    i_014    tia_h_in_001_019+    119396.17708026717
Rh001_014_019-    i_014    tia_h_in_001_019-    76311.2289124319
Rh001_015_019+    i_015    tia_h_in_001_019+    120359.67015579385
Rh001_015_019-    i_015    tia_h_in_001_019-    66195.56040027601
Rh001_016_019+    i_016    tia_h_in_001_019+    67544.14427359092
Rh001_016_019-    i_016    tia_h_in_001_019-    119302.88344931396
Rh001_017_019+    i_017    tia_h_in_001_019+    31993.477556668502
Rh001_017_019-    i_017    tia_h_in_001_019-    120000
Rh001_018_019+    i_018    tia_h_in_001_019+    32925.286825495044
Rh001_018_019-    i_018    tia_h_in_001_019-    118481.24977169957
Rh001_019_019+    i_019    tia_h_in_001_019+    85263.20173375023
Rh001_019_019-    i_019    tia_h_in_001_019-    119528.87386114206
Rh001_020_019+    i_020    tia_h_in_001_019+    102018.34278199782
Rh001_020_019-    i_020    tia_h_in_001_019-    118446.50566967452
Rh001_021_019+    i_021    tia_h_in_001_019+    118720.58834404727
Rh001_021_019-    i_021    tia_h_in_001_019-    56167.82400497889
Rh001_022_019+    i_022    tia_h_in_001_019+    121065.81064044456
Rh001_022_019-    i_022    tia_h_in_001_019-    68248.69189580943
Rh001_023_019+    i_023    tia_h_in_001_019+    102728.45404514021
Rh001_023_019-    i_023    tia_h_in_001_019-    120786.19633922196
Rh001_024_019+    i_024    tia_h_in_001_019+    70007.51686089796
Rh001_024_019-    i_024    tia_h_in_001_019-    119001.76934935813
Rh001_025_019+    i_025    tia_h_in_001_019+    36115.34485504362
Rh001_025_019-    i_025    tia_h_in_001_019-    120678.98870543447
Rh001_026_019+    i_026    tia_h_in_001_019+    5000
Rh001_026_019-    i_026    tia_h_in_001_019-    5000
Rh001_027_019+    i_027    tia_h_in_001_019+    119176.5264596186
Rh001_027_019-    i_027    tia_h_in_001_019-    49466.77186536819
Rh001_028_019+    i_028    tia_h_in_001_019+    120804.48409671675
Rh001_028_019-    i_028    tia_h_in_001_019-    80402.71255518546
Rh001_029_019+    i_029    tia_h_in_001_019+    121345.37428998714
Rh001_029_019-    i_029    tia_h_in_001_019-    51882.37996473427
Rh001_030_019+    i_030    tia_h_in_001_019+    120831.86826909952
Rh001_030_019-    i_030    tia_h_in_001_019-    50544.362562484115
Rh001_031_019+    i_031    tia_h_in_001_019+    62543.38380431629
Rh001_031_019-    i_031    tia_h_in_001_019-    121790.99948080232
Rh001_032_019+    i_032    tia_h_in_001_019+    55801.4033442031
Rh001_032_019-    i_032    tia_h_in_001_019-    119456.25926863546
Rh001_033_019+    i_033    tia_h_in_001_019+    64229.197075206794
Rh001_033_019-    i_033    tia_h_in_001_019-    120645.53960491886
Rh001_034_019+    i_034    tia_h_in_001_019+    82559.84951723776
Rh001_034_019-    i_034    tia_h_in_001_019-    121581.1705614735
Rh001_035_019+    i_035    tia_h_in_001_019+    118644.1082149823
Rh001_035_019-    i_035    tia_h_in_001_019-    61841.3218070022
Rh001_036_019+    i_036    tia_h_in_001_019+    120852.355778058
Rh001_036_019-    i_036    tia_h_in_001_019-    54106.09650412362
Rh001_037_019+    i_037    tia_h_in_001_019+    5000
Rh001_037_019-    i_037    tia_h_in_001_019-    46121.22161945601
Rh001_038_019+    i_038    tia_h_in_001_019+    64213.19031885574
Rh001_038_019-    i_038    tia_h_in_001_019-    119540.59450009049
Rh001_039_019+    i_039    tia_h_in_001_019+    120964.47811993635
Rh001_039_019-    i_039    tia_h_in_001_019-    115510.26576243578
Rh001_040_019+    i_040    tia_h_in_001_019+    43962.1127331437
Rh001_040_019-    i_040    tia_h_in_001_019-    120101.050666841
Rh001_041_019+    i_041    tia_h_in_001_019+    120903.97166667238
Rh001_041_019-    i_041    tia_h_in_001_019-    54451.115140709255
Rh001_042_019+    i_042    tia_h_in_001_019+    120370.21529235509
Rh001_042_019-    i_042    tia_h_in_001_019-    120000
Rh001_043_019+    i_043    tia_h_in_001_019+    122087.92243013937
Rh001_043_019-    i_043    tia_h_in_001_019-    44130.418885226485
Rh001_044_019+    i_044    tia_h_in_001_019+    119621.5390783061
Rh001_044_019-    i_044    tia_h_in_001_019-    117954.61506785225
Rh001_045_019+    i_045    tia_h_in_001_019+    5000
Rh001_045_019-    i_045    tia_h_in_001_019-    120393.37439979428
Rh001_046_019+    i_046    tia_h_in_001_019+    36659.10918421978
Rh001_046_019-    i_046    tia_h_in_001_019-    120164.04650164477
Rh001_047_019+    i_047    tia_h_in_001_019+    65377.683544460844
Rh001_047_019-    i_047    tia_h_in_001_019-    119827.32720019699
Rh001_048_019+    i_048    tia_h_in_001_019+    67730.60016392764
Rh001_048_019-    i_048    tia_h_in_001_019-    119805.84353947877
Rh001_049_019+    i_049    tia_h_in_001_019+    119693.93329430801
Rh001_049_019-    i_049    tia_h_in_001_019-    51926.56327978594
Rh001_050_019+    i_050    tia_h_in_001_019+    118184.10421238594
Rh001_050_019-    i_050    tia_h_in_001_019-    42568.571148815965
Rh001_051_019+    i_051    tia_h_in_001_019+    119296.78608407317
Rh001_051_019-    i_051    tia_h_in_001_019-    42773.901764689275
Rh001_052_019+    i_052    tia_h_in_001_019+    114966.86292105899
Rh001_052_019-    i_052    tia_h_in_001_019-    119029.48814404392
Rh001_053_019+    i_053    tia_h_in_001_019+    119914.01452539918
Rh001_053_019-    i_053    tia_h_in_001_019-    113937.531019822
Rh001_054_019+    i_054    tia_h_in_001_019+    43017.936197476934
Rh001_054_019-    i_054    tia_h_in_001_019-    119507.37519385586
Rh001_055_019+    i_055    tia_h_in_001_019+    32329.647951539835
Rh001_055_019-    i_055    tia_h_in_001_019-    119769.9978037549
Rh001_056_019+    i_056    tia_h_in_001_019+    117247.75400699688
Rh001_056_019-    i_056    tia_h_in_001_019-    119333.10440013462
Rh001_057_019+    i_057    tia_h_in_001_019+    120846.29851835736
Rh001_057_019-    i_057    tia_h_in_001_019-    21142.732144711455
Rh001_058_019+    i_058    tia_h_in_001_019+    118949.96818650466
Rh001_058_019-    i_058    tia_h_in_001_019-    41739.722460222605
Rh001_059_019+    i_059    tia_h_in_001_019+    118731.03568939018
Rh001_059_019-    i_059    tia_h_in_001_019-    89290.12541750398
Rh001_060_019+    i_060    tia_h_in_001_019+    26275.23836362052
Rh001_060_019-    i_060    tia_h_in_001_019-    122117.03986870003
Rh001_061_019+    i_061    tia_h_in_001_019+    17193.27772117594
Rh001_061_019-    i_061    tia_h_in_001_019-    118400.6299423771
Rh001_062_019+    i_062    tia_h_in_001_019+    29773.99200490035
Rh001_062_019-    i_062    tia_h_in_001_019-    119147.45375745077
Rh001_063_019+    i_063    tia_h_in_001_019+    118858.63362406654
Rh001_063_019-    i_063    tia_h_in_001_019-    51791.128542526305
Rh001_064_019+    i_064    tia_h_in_001_019+    119211.38294002232
Rh001_064_019-    i_064    tia_h_in_001_019-    120000

* Neuron 20
Rh001_001_020+    i_001    tia_h_in_001_020+    119398.90413965924
Rh001_001_020-    i_001    tia_h_in_001_020-    45928.751897946015
Rh001_002_020+    i_002    tia_h_in_001_020+    120436.16709285467
Rh001_002_020-    i_002    tia_h_in_001_020-    39802.7313216204
Rh001_003_020+    i_003    tia_h_in_001_020+    120618.05858312843
Rh001_003_020-    i_003    tia_h_in_001_020-    33123.52607449434
Rh001_004_020+    i_004    tia_h_in_001_020+    5000
Rh001_004_020-    i_004    tia_h_in_001_020-    120366.49348081727
Rh001_005_020+    i_005    tia_h_in_001_020+    119597.90028935569
Rh001_005_020-    i_005    tia_h_in_001_020-    5000
Rh001_006_020+    i_006    tia_h_in_001_020+    59690.28296077333
Rh001_006_020-    i_006    tia_h_in_001_020-    120000
Rh001_007_020+    i_007    tia_h_in_001_020+    40681.60055628521
Rh001_007_020-    i_007    tia_h_in_001_020-    119248.45651024458
Rh001_008_020+    i_008    tia_h_in_001_020+    41266.74412090154
Rh001_008_020-    i_008    tia_h_in_001_020-    119843.7927918303
Rh001_009_020+    i_009    tia_h_in_001_020+    110263.6586752628
Rh001_009_020-    i_009    tia_h_in_001_020-    118182.241864025
Rh001_010_020+    i_010    tia_h_in_001_020+    119450.87056903719
Rh001_010_020-    i_010    tia_h_in_001_020-    25305.127748655766
Rh001_011_020+    i_011    tia_h_in_001_020+    31865.03657631271
Rh001_011_020-    i_011    tia_h_in_001_020-    120000
Rh001_012_020+    i_012    tia_h_in_001_020+    39817.6426071136
Rh001_012_020-    i_012    tia_h_in_001_020-    120595.82519122383
Rh001_013_020+    i_013    tia_h_in_001_020+    122567.41117944074
Rh001_013_020-    i_013    tia_h_in_001_020-    87308.70461682565
Rh001_014_020+    i_014    tia_h_in_001_020+    40036.70457668181
Rh001_014_020-    i_014    tia_h_in_001_020-    120933.55888725712
Rh001_015_020+    i_015    tia_h_in_001_020+    79808.5622343688
Rh001_015_020-    i_015    tia_h_in_001_020-    119216.69240057103
Rh001_016_020+    i_016    tia_h_in_001_020+    5000
Rh001_016_020-    i_016    tia_h_in_001_020-    121380.79955073305
Rh001_017_020+    i_017    tia_h_in_001_020+    120543.45946669672
Rh001_017_020-    i_017    tia_h_in_001_020-    32882.96011054367
Rh001_018_020+    i_018    tia_h_in_001_020+    74497.4001934948
Rh001_018_020-    i_018    tia_h_in_001_020-    117605.98327633984
Rh001_019_020+    i_019    tia_h_in_001_020+    61222.3878902236
Rh001_019_020-    i_019    tia_h_in_001_020-    121154.13348833131
Rh001_020_020+    i_020    tia_h_in_001_020+    55923.406256254
Rh001_020_020-    i_020    tia_h_in_001_020-    120173.81418307949
Rh001_021_020+    i_021    tia_h_in_001_020+    119447.84443479858
Rh001_021_020-    i_021    tia_h_in_001_020-    90417.14453288255
Rh001_022_020+    i_022    tia_h_in_001_020+    121333.7905049688
Rh001_022_020-    i_022    tia_h_in_001_020-    86294.03921512743
Rh001_023_020+    i_023    tia_h_in_001_020+    85201.34762554058
Rh001_023_020-    i_023    tia_h_in_001_020-    121756.628164513
Rh001_024_020+    i_024    tia_h_in_001_020+    42708.55045800013
Rh001_024_020-    i_024    tia_h_in_001_020-    120451.20889530549
Rh001_025_020+    i_025    tia_h_in_001_020+    107604.06770357325
Rh001_025_020-    i_025    tia_h_in_001_020-    5000
Rh001_026_020+    i_026    tia_h_in_001_020+    95894.767104254
Rh001_026_020-    i_026    tia_h_in_001_020-    120920.01128271478
Rh001_027_020+    i_027    tia_h_in_001_020+    119972.39678982693
Rh001_027_020-    i_027    tia_h_in_001_020-    76483.91030667654
Rh001_028_020+    i_028    tia_h_in_001_020+    120344.15112943946
Rh001_028_020-    i_028    tia_h_in_001_020-    36084.34106272476
Rh001_029_020+    i_029    tia_h_in_001_020+    118575.65649849064
Rh001_029_020-    i_029    tia_h_in_001_020-    53091.93220334666
Rh001_030_020+    i_030    tia_h_in_001_020+    119594.81608041115
Rh001_030_020-    i_030    tia_h_in_001_020-    67369.82783797165
Rh001_031_020+    i_031    tia_h_in_001_020+    119709.56907035763
Rh001_031_020-    i_031    tia_h_in_001_020-    62417.34895502716
Rh001_032_020+    i_032    tia_h_in_001_020+    105698.67320223396
Rh001_032_020-    i_032    tia_h_in_001_020-    120409.24524997178
Rh001_033_020+    i_033    tia_h_in_001_020+    91163.65369130624
Rh001_033_020-    i_033    tia_h_in_001_020-    120764.41391303796
Rh001_034_020+    i_034    tia_h_in_001_020+    121772.90037965593
Rh001_034_020-    i_034    tia_h_in_001_020-    84121.13824587267
Rh001_035_020+    i_035    tia_h_in_001_020+    120000
Rh001_035_020-    i_035    tia_h_in_001_020-    119139.94226204249
Rh001_036_020+    i_036    tia_h_in_001_020+    120245.87258573835
Rh001_036_020-    i_036    tia_h_in_001_020-    64082.86085825511
Rh001_037_020+    i_037    tia_h_in_001_020+    119632.64424880216
Rh001_037_020-    i_037    tia_h_in_001_020-    47117.32034795498
Rh001_038_020+    i_038    tia_h_in_001_020+    80103.00586828806
Rh001_038_020-    i_038    tia_h_in_001_020-    121133.01479060666
Rh001_039_020+    i_039    tia_h_in_001_020+    68607.29528699984
Rh001_039_020-    i_039    tia_h_in_001_020-    119018.73527521155
Rh001_040_020+    i_040    tia_h_in_001_020+    121816.60101984435
Rh001_040_020-    i_040    tia_h_in_001_020-    51218.20169084074
Rh001_041_020+    i_041    tia_h_in_001_020+    93373.26038219711
Rh001_041_020-    i_041    tia_h_in_001_020-    5000
Rh001_042_020+    i_042    tia_h_in_001_020+    5000
Rh001_042_020-    i_042    tia_h_in_001_020-    119614.16375240198
Rh001_043_020+    i_043    tia_h_in_001_020+    120106.97811470627
Rh001_043_020-    i_043    tia_h_in_001_020-    37047.427574109686
Rh001_044_020+    i_044    tia_h_in_001_020+    119743.9028007835
Rh001_044_020-    i_044    tia_h_in_001_020-    47542.99055017713
Rh001_045_020+    i_045    tia_h_in_001_020+    120000
Rh001_045_020-    i_045    tia_h_in_001_020-    121152.40439494014
Rh001_046_020+    i_046    tia_h_in_001_020+    50679.2155709423
Rh001_046_020-    i_046    tia_h_in_001_020-    121384.21849960246
Rh001_047_020+    i_047    tia_h_in_001_020+    54016.555023376975
Rh001_047_020-    i_047    tia_h_in_001_020-    118944.1310048093
Rh001_048_020+    i_048    tia_h_in_001_020+    118521.40261954577
Rh001_048_020-    i_048    tia_h_in_001_020-    104527.0005774943
Rh001_049_020+    i_049    tia_h_in_001_020+    52153.17143998118
Rh001_049_020-    i_049    tia_h_in_001_020-    5000
Rh001_050_020+    i_050    tia_h_in_001_020+    5000
Rh001_050_020-    i_050    tia_h_in_001_020-    118870.48764541157
Rh001_051_020+    i_051    tia_h_in_001_020+    40508.89214212851
Rh001_051_020-    i_051    tia_h_in_001_020-    120642.91395079435
Rh001_052_020+    i_052    tia_h_in_001_020+    56511.62168987871
Rh001_052_020-    i_052    tia_h_in_001_020-    119764.82802251617
Rh001_053_020+    i_053    tia_h_in_001_020+    92073.83685036091
Rh001_053_020-    i_053    tia_h_in_001_020-    120000
Rh001_054_020+    i_054    tia_h_in_001_020+    55196.97430950747
Rh001_054_020-    i_054    tia_h_in_001_020-    120031.96221618557
Rh001_055_020+    i_055    tia_h_in_001_020+    119943.80564184827
Rh001_055_020-    i_055    tia_h_in_001_020-    31156.065686812588
Rh001_056_020+    i_056    tia_h_in_001_020+    121202.29255065005
Rh001_056_020-    i_056    tia_h_in_001_020-    77112.27220738167
Rh001_057_020+    i_057    tia_h_in_001_020+    45332.93198589533
Rh001_057_020-    i_057    tia_h_in_001_020-    120000
Rh001_058_020+    i_058    tia_h_in_001_020+    63787.90250508852
Rh001_058_020-    i_058    tia_h_in_001_020-    120321.14497222142
Rh001_059_020+    i_059    tia_h_in_001_020+    37480.46065009718
Rh001_059_020-    i_059    tia_h_in_001_020-    121664.18822598459
Rh001_060_020+    i_060    tia_h_in_001_020+    98807.03258710178
Rh001_060_020-    i_060    tia_h_in_001_020-    120613.04940660493
Rh001_061_020+    i_061    tia_h_in_001_020+    110745.95175458789
Rh001_061_020-    i_061    tia_h_in_001_020-    120000
Rh001_062_020+    i_062    tia_h_in_001_020+    119846.97570628974
Rh001_062_020-    i_062    tia_h_in_001_020-    35593.58022859293
Rh001_063_020+    i_063    tia_h_in_001_020+    119863.69520909767
Rh001_063_020-    i_063    tia_h_in_001_020-    26561.406139952585
Rh001_064_020+    i_064    tia_h_in_001_020+    120278.43215102854
Rh001_064_020-    i_064    tia_h_in_001_020-    120000

* ----- Bias
    
        
Rb_h001_001+    b_001    tia_h_in_001_001+    120627.1642634071
Rb_h001_001-    b_001    tia_h_in_001_001-    120000
Rb_h001_002+    b_001    tia_h_in_001_002+    28980.64763141459
Rb_h001_002-    b_001    tia_h_in_001_002-    120435.73315254063
Rb_h001_003+    b_001    tia_h_in_001_003+    120367.10851147871
Rb_h001_003-    b_001    tia_h_in_001_003-    16016.173678873034
Rb_h001_004+    b_001    tia_h_in_001_004+    120488.84074450962
Rb_h001_004-    b_001    tia_h_in_001_004-    54091.01002265623
Rb_h001_005+    b_001    tia_h_in_001_005+    5000
Rb_h001_005-    b_001    tia_h_in_001_005-    120638.11515493115
Rb_h001_006+    b_001    tia_h_in_001_006+    82981.47977793262
Rb_h001_006-    b_001    tia_h_in_001_006-    119350.76893994444
Rb_h001_007+    b_001    tia_h_in_001_007+    47010.515167273385
Rb_h001_007-    b_001    tia_h_in_001_007-    120747.8414145181
Rb_h001_008+    b_001    tia_h_in_001_008+    43240.013507893884
Rb_h001_008-    b_001    tia_h_in_001_008-    119168.06674257849
Rb_h001_009+    b_001    tia_h_in_001_009+    31982.441119856587
Rb_h001_009-    b_001    tia_h_in_001_009-    121303.60646207984
Rb_h001_010+    b_001    tia_h_in_001_010+    120882.17736444659
Rb_h001_010-    b_001    tia_h_in_001_010-    81629.19162800473
Rb_h001_011+    b_001    tia_h_in_001_011+    35683.55385848612
Rb_h001_011-    b_001    tia_h_in_001_011-    120182.25375768416
Rb_h001_012+    b_001    tia_h_in_001_012+    26375.664431244564
Rb_h001_012-    b_001    tia_h_in_001_012-    120336.19207207374
Rb_h001_013+    b_001    tia_h_in_001_013+    61128.78613467687
Rb_h001_013-    b_001    tia_h_in_001_013-    120607.56585862239
Rb_h001_014+    b_001    tia_h_in_001_014+    120869.71017527606
Rb_h001_014-    b_001    tia_h_in_001_014-    54838.43522597561
Rb_h001_015+    b_001    tia_h_in_001_015+    120000
Rb_h001_015-    b_001    tia_h_in_001_015-    120563.96816122452
Rb_h001_016+    b_001    tia_h_in_001_016+    120107.09215569988
Rb_h001_016-    b_001    tia_h_in_001_016-    34335.10161759296
Rb_h001_017+    b_001    tia_h_in_001_017+    120738.52513062558
Rb_h001_017-    b_001    tia_h_in_001_017-    47803.13952471517
Rb_h001_018+    b_001    tia_h_in_001_018+    5000
Rb_h001_018-    b_001    tia_h_in_001_018-    121124.26020110332
Rb_h001_019+    b_001    tia_h_in_001_019+    119498.16142786323
Rb_h001_019-    b_001    tia_h_in_001_019-    15825.633712116887
Rb_h001_020+    b_001    tia_h_in_001_020+    28819.304212178824
Rb_h001_020-    b_001    tia_h_in_001_020-    121405.58130045343

* ----- Weights
* Layer 002

* Neuron 1
Rh002_001_001+    hidden_activ_out_h001_001    tia_h_in_002_001+    5000
Rh002_001_001-    hidden_activ_out_h001_001    tia_h_in_002_001-    7356.515850321617
Rh002_002_001+    hidden_activ_out_h001_002    tia_h_in_002_001+    5000
Rh002_002_001-    hidden_activ_out_h001_002    tia_h_in_002_001-    120297.21238648427
Rh002_003_001+    hidden_activ_out_h001_003    tia_h_in_002_001+    119051.77541642915
Rh002_003_001-    hidden_activ_out_h001_003    tia_h_in_002_001-    7322.286566428803
Rh002_004_001+    hidden_activ_out_h001_004    tia_h_in_002_001+    5000
Rh002_004_001-    hidden_activ_out_h001_004    tia_h_in_002_001-    45497.72992256005
Rh002_005_001+    hidden_activ_out_h001_005    tia_h_in_002_001+    6042.024578583226
Rh002_005_001-    hidden_activ_out_h001_005    tia_h_in_002_001-    121681.70512346842
Rh002_006_001+    hidden_activ_out_h001_006    tia_h_in_002_001+    120784.41367394988
Rh002_006_001-    hidden_activ_out_h001_006    tia_h_in_002_001-    112216.69190444781
Rh002_007_001+    hidden_activ_out_h001_007    tia_h_in_002_001+    26602.844191391894
Rh002_007_001-    hidden_activ_out_h001_007    tia_h_in_002_001-    119889.6256745405
Rh002_008_001+    hidden_activ_out_h001_008    tia_h_in_002_001+    6488.135254704738
Rh002_008_001-    hidden_activ_out_h001_008    tia_h_in_002_001-    121123.0199287729
Rh002_009_001+    hidden_activ_out_h001_009    tia_h_in_002_001+    19824.301399182732
Rh002_009_001-    hidden_activ_out_h001_009    tia_h_in_002_001-    119645.11154887384
Rh002_010_001+    hidden_activ_out_h001_010    tia_h_in_002_001+    121396.66398909784
Rh002_010_001-    hidden_activ_out_h001_010    tia_h_in_002_001-    79711.16467831444
Rh002_011_001+    hidden_activ_out_h001_011    tia_h_in_002_001+    11695.769264885737
Rh002_011_001-    hidden_activ_out_h001_011    tia_h_in_002_001-    119088.72484680454
Rh002_012_001+    hidden_activ_out_h001_012    tia_h_in_002_001+    120892.63527838663
Rh002_012_001-    hidden_activ_out_h001_012    tia_h_in_002_001-    5000
Rh002_013_001+    hidden_activ_out_h001_013    tia_h_in_002_001+    11955.453640873062
Rh002_013_001-    hidden_activ_out_h001_013    tia_h_in_002_001-    120689.65242807804
Rh002_014_001+    hidden_activ_out_h001_014    tia_h_in_002_001+    122914.06367642427
Rh002_014_001-    hidden_activ_out_h001_014    tia_h_in_002_001-    118312.76417560023
Rh002_015_001+    hidden_activ_out_h001_015    tia_h_in_002_001+    119725.6091972224
Rh002_015_001-    hidden_activ_out_h001_015    tia_h_in_002_001-    120000
Rh002_016_001+    hidden_activ_out_h001_016    tia_h_in_002_001+    120230.86524181587
Rh002_016_001-    hidden_activ_out_h001_016    tia_h_in_002_001-    8598.703664192384
Rh002_017_001+    hidden_activ_out_h001_017    tia_h_in_002_001+    121085.37972738099
Rh002_017_001-    hidden_activ_out_h001_017    tia_h_in_002_001-    7739.397244461697
Rh002_018_001+    hidden_activ_out_h001_018    tia_h_in_002_001+    29966.169739297795
Rh002_018_001-    hidden_activ_out_h001_018    tia_h_in_002_001-    119522.44742760435
Rh002_019_001+    hidden_activ_out_h001_019    tia_h_in_002_001+    120666.42785947006
Rh002_019_001-    hidden_activ_out_h001_019    tia_h_in_002_001-    6602.951624177698
Rh002_020_001+    hidden_activ_out_h001_020    tia_h_in_002_001+    120962.69945800917
Rh002_020_001-    hidden_activ_out_h001_020    tia_h_in_002_001-    120000

* Neuron 2
Rh002_001_002+    hidden_activ_out_h001_001    tia_h_in_002_002+    119996.87753430833
Rh002_001_002-    hidden_activ_out_h001_001    tia_h_in_002_002-    29092.34292985449
Rh002_002_002+    hidden_activ_out_h001_002    tia_h_in_002_002+    119894.42989342174
Rh002_002_002-    hidden_activ_out_h001_002    tia_h_in_002_002-    120000
Rh002_003_002+    hidden_activ_out_h001_003    tia_h_in_002_002+    18231.94624464673
Rh002_003_002-    hidden_activ_out_h001_003    tia_h_in_002_002-    120668.46109653433
Rh002_004_002+    hidden_activ_out_h001_004    tia_h_in_002_002+    41355.04044200833
Rh002_004_002-    hidden_activ_out_h001_004    tia_h_in_002_002-    120793.68898810036
Rh002_005_002+    hidden_activ_out_h001_005    tia_h_in_002_002+    120321.82131367568
Rh002_005_002-    hidden_activ_out_h001_005    tia_h_in_002_002-    10569.172208677926
Rh002_006_002+    hidden_activ_out_h001_006    tia_h_in_002_002+    66893.62996130773
Rh002_006_002-    hidden_activ_out_h001_006    tia_h_in_002_002-    118156.76356952715
Rh002_007_002+    hidden_activ_out_h001_007    tia_h_in_002_002+    121243.8207497502
Rh002_007_002-    hidden_activ_out_h001_007    tia_h_in_002_002-    9153.373623583195
Rh002_008_002+    hidden_activ_out_h001_008    tia_h_in_002_002+    121126.13821104044
Rh002_008_002-    hidden_activ_out_h001_008    tia_h_in_002_002-    9313.473820215986
Rh002_009_002+    hidden_activ_out_h001_009    tia_h_in_002_002+    119590.15473123326
Rh002_009_002-    hidden_activ_out_h001_009    tia_h_in_002_002-    9285.968857386722
Rh002_010_002+    hidden_activ_out_h001_010    tia_h_in_002_002+    44691.347923364854
Rh002_010_002-    hidden_activ_out_h001_010    tia_h_in_002_002-    117451.15018812541
Rh002_011_002+    hidden_activ_out_h001_011    tia_h_in_002_002+    122350.55161702592
Rh002_011_002-    hidden_activ_out_h001_011    tia_h_in_002_002-    8781.717141372728
Rh002_012_002+    hidden_activ_out_h001_012    tia_h_in_002_002+    120899.54454282622
Rh002_012_002-    hidden_activ_out_h001_012    tia_h_in_002_002-    16767.286723921414
Rh002_013_002+    hidden_activ_out_h001_013    tia_h_in_002_002+    120212.06558499018
Rh002_013_002-    hidden_activ_out_h001_013    tia_h_in_002_002-    7954.7622380744815
Rh002_014_002+    hidden_activ_out_h001_014    tia_h_in_002_002+    120203.59853838774
Rh002_014_002-    hidden_activ_out_h001_014    tia_h_in_002_002-    81075.36510947357
Rh002_015_002+    hidden_activ_out_h001_015    tia_h_in_002_002+    37869.27648294926
Rh002_015_002-    hidden_activ_out_h001_015    tia_h_in_002_002-    119258.3040364719
Rh002_016_002+    hidden_activ_out_h001_016    tia_h_in_002_002+    119498.02180790043
Rh002_016_002-    hidden_activ_out_h001_016    tia_h_in_002_002-    120000
Rh002_017_002+    hidden_activ_out_h001_017    tia_h_in_002_002+    94242.44196138643
Rh002_017_002-    hidden_activ_out_h001_017    tia_h_in_002_002-    120974.53013285412
Rh002_018_002+    hidden_activ_out_h001_018    tia_h_in_002_002+    121183.7508734986
Rh002_018_002-    hidden_activ_out_h001_018    tia_h_in_002_002-    7761.366806990562
Rh002_019_002+    hidden_activ_out_h001_019    tia_h_in_002_002+    16447.005495755555
Rh002_019_002-    hidden_activ_out_h001_019    tia_h_in_002_002-    119749.93411576588
Rh002_020_002+    hidden_activ_out_h001_020    tia_h_in_002_002+    117967.4215273276
Rh002_020_002-    hidden_activ_out_h001_020    tia_h_in_002_002-    10707.4804130226

* Neuron 3
Rh002_001_003+    hidden_activ_out_h001_001    tia_h_in_002_003+    18563.057585824325
Rh002_001_003-    hidden_activ_out_h001_001    tia_h_in_002_003-    120077.01373965283
Rh002_002_003+    hidden_activ_out_h001_002    tia_h_in_002_003+    120447.21491176852
Rh002_002_003-    hidden_activ_out_h001_002    tia_h_in_002_003-    7392.554535824334
Rh002_003_003+    hidden_activ_out_h001_003    tia_h_in_002_003+    33914.86797392436
Rh002_003_003-    hidden_activ_out_h001_003    tia_h_in_002_003-    119607.86366613742
Rh002_004_003+    hidden_activ_out_h001_004    tia_h_in_002_003+    69067.96467186067
Rh002_004_003-    hidden_activ_out_h001_004    tia_h_in_002_003-    121030.53919969186
Rh002_005_003+    hidden_activ_out_h001_005    tia_h_in_002_003+    119905.79698192317
Rh002_005_003-    hidden_activ_out_h001_005    tia_h_in_002_003-    13434.782503098659
Rh002_006_003+    hidden_activ_out_h001_006    tia_h_in_002_003+    121714.61153319848
Rh002_006_003-    hidden_activ_out_h001_006    tia_h_in_002_003-    85884.27979448024
Rh002_007_003+    hidden_activ_out_h001_007    tia_h_in_002_003+    120730.3194387346
Rh002_007_003-    hidden_activ_out_h001_007    tia_h_in_002_003-    16214.897004693212
Rh002_008_003+    hidden_activ_out_h001_008    tia_h_in_002_003+    120047.55652498697
Rh002_008_003-    hidden_activ_out_h001_008    tia_h_in_002_003-    19323.667983955
Rh002_009_003+    hidden_activ_out_h001_009    tia_h_in_002_003+    122188.54087495533
Rh002_009_003-    hidden_activ_out_h001_009    tia_h_in_002_003-    10687.406738258172
Rh002_010_003+    hidden_activ_out_h001_010    tia_h_in_002_003+    106355.78485084457
Rh002_010_003-    hidden_activ_out_h001_010    tia_h_in_002_003-    5000
Rh002_011_003+    hidden_activ_out_h001_011    tia_h_in_002_003+    121253.51299049146
Rh002_011_003-    hidden_activ_out_h001_011    tia_h_in_002_003-    11498.210848736331
Rh002_012_003+    hidden_activ_out_h001_012    tia_h_in_002_003+    120000
Rh002_012_003-    hidden_activ_out_h001_012    tia_h_in_002_003-    21676.308723119524
Rh002_013_003+    hidden_activ_out_h001_013    tia_h_in_002_003+    119530.82126428408
Rh002_013_003-    hidden_activ_out_h001_013    tia_h_in_002_003-    10595.624690937535
Rh002_014_003+    hidden_activ_out_h001_014    tia_h_in_002_003+    48448.43192233514
Rh002_014_003-    hidden_activ_out_h001_014    tia_h_in_002_003-    119329.97299168208
Rh002_015_003+    hidden_activ_out_h001_015    tia_h_in_002_003+    96968.02517164945
Rh002_015_003-    hidden_activ_out_h001_015    tia_h_in_002_003-    120661.38839162397
Rh002_016_003+    hidden_activ_out_h001_016    tia_h_in_002_003+    19911.763119238058
Rh002_016_003-    hidden_activ_out_h001_016    tia_h_in_002_003-    119638.1338048662
Rh002_017_003+    hidden_activ_out_h001_017    tia_h_in_002_003+    120202.91816649678
Rh002_017_003-    hidden_activ_out_h001_017    tia_h_in_002_003-    18245.224267815654
Rh002_018_003+    hidden_activ_out_h001_018    tia_h_in_002_003+    119449.33103610884
Rh002_018_003-    hidden_activ_out_h001_018    tia_h_in_002_003-    17592.662389908317
Rh002_019_003+    hidden_activ_out_h001_019    tia_h_in_002_003+    43306.04441432542
Rh002_019_003-    hidden_activ_out_h001_019    tia_h_in_002_003-    122119.92317286413
Rh002_020_003+    hidden_activ_out_h001_020    tia_h_in_002_003+    119916.29303768373
Rh002_020_003-    hidden_activ_out_h001_020    tia_h_in_002_003-    32990.837293328535

* Neuron 4
Rh002_001_004+    hidden_activ_out_h001_001    tia_h_in_002_004+    120000
Rh002_001_004-    hidden_activ_out_h001_001    tia_h_in_002_004-    120704.03938794282
Rh002_002_004+    hidden_activ_out_h001_002    tia_h_in_002_004+    120096.15687356405
Rh002_002_004-    hidden_activ_out_h001_002    tia_h_in_002_004-    20585.764215792922
Rh002_003_004+    hidden_activ_out_h001_003    tia_h_in_002_004+    22754.188383963654
Rh002_003_004-    hidden_activ_out_h001_003    tia_h_in_002_004-    120136.42484604713
Rh002_004_004+    hidden_activ_out_h001_004    tia_h_in_002_004+    119705.41663202927
Rh002_004_004-    hidden_activ_out_h001_004    tia_h_in_002_004-    44510.08716253386
Rh002_005_004+    hidden_activ_out_h001_005    tia_h_in_002_004+    120336.48111803898
Rh002_005_004-    hidden_activ_out_h001_005    tia_h_in_002_004-    16317.910272310228
Rh002_006_004+    hidden_activ_out_h001_006    tia_h_in_002_004+    5000
Rh002_006_004-    hidden_activ_out_h001_006    tia_h_in_002_004-    118993.6616662024
Rh002_007_004+    hidden_activ_out_h001_007    tia_h_in_002_004+    118282.01343527742
Rh002_007_004-    hidden_activ_out_h001_007    tia_h_in_002_004-    26626.554450249303
Rh002_008_004+    hidden_activ_out_h001_008    tia_h_in_002_004+    120755.08501867761
Rh002_008_004-    hidden_activ_out_h001_008    tia_h_in_002_004-    120000
Rh002_009_004+    hidden_activ_out_h001_009    tia_h_in_002_004+    122188.93829217106
Rh002_009_004-    hidden_activ_out_h001_009    tia_h_in_002_004-    60341.93084099196
Rh002_010_004+    hidden_activ_out_h001_010    tia_h_in_002_004+    120445.6613740111
Rh002_010_004-    hidden_activ_out_h001_010    tia_h_in_002_004-    38561.096214943755
Rh002_011_004+    hidden_activ_out_h001_011    tia_h_in_002_004+    121622.98886939227
Rh002_011_004-    hidden_activ_out_h001_011    tia_h_in_002_004-    26533.960353768656
Rh002_012_004+    hidden_activ_out_h001_012    tia_h_in_002_004+    119413.04497841565
Rh002_012_004-    hidden_activ_out_h001_012    tia_h_in_002_004-    5000
Rh002_013_004+    hidden_activ_out_h001_013    tia_h_in_002_004+    120312.22875610962
Rh002_013_004-    hidden_activ_out_h001_013    tia_h_in_002_004-    32159.40417691629
Rh002_014_004+    hidden_activ_out_h001_014    tia_h_in_002_004+    120330.2747048637
Rh002_014_004-    hidden_activ_out_h001_014    tia_h_in_002_004-    75121.70673781745
Rh002_015_004+    hidden_activ_out_h001_015    tia_h_in_002_004+    45173.50729806501
Rh002_015_004-    hidden_activ_out_h001_015    tia_h_in_002_004-    120910.2199723631
Rh002_016_004+    hidden_activ_out_h001_016    tia_h_in_002_004+    13049.520979373541
Rh002_016_004-    hidden_activ_out_h001_016    tia_h_in_002_004-    120057.67425529876
Rh002_017_004+    hidden_activ_out_h001_017    tia_h_in_002_004+    5000
Rh002_017_004-    hidden_activ_out_h001_017    tia_h_in_002_004-    120363.5789053314
Rh002_018_004+    hidden_activ_out_h001_018    tia_h_in_002_004+    120000
Rh002_018_004-    hidden_activ_out_h001_018    tia_h_in_002_004-    69676.7983837342
Rh002_019_004+    hidden_activ_out_h001_019    tia_h_in_002_004+    15402.126613566788
Rh002_019_004-    hidden_activ_out_h001_019    tia_h_in_002_004-    119099.12347225899
Rh002_020_004+    hidden_activ_out_h001_020    tia_h_in_002_004+    119060.25381253492
Rh002_020_004-    hidden_activ_out_h001_020    tia_h_in_002_004-    94829.87885636455

* Neuron 5
Rh002_001_005+    hidden_activ_out_h001_001    tia_h_in_002_005+    15774.50964345318
Rh002_001_005-    hidden_activ_out_h001_001    tia_h_in_002_005-    119579.49494957857
Rh002_002_005+    hidden_activ_out_h001_002    tia_h_in_002_005+    119870.97454997581
Rh002_002_005-    hidden_activ_out_h001_002    tia_h_in_002_005-    19623.1554399893
Rh002_003_005+    hidden_activ_out_h001_003    tia_h_in_002_005+    28525.060131899278
Rh002_003_005-    hidden_activ_out_h001_003    tia_h_in_002_005-    119338.09341471083
Rh002_004_005+    hidden_activ_out_h001_004    tia_h_in_002_005+    77279.7500550574
Rh002_004_005-    hidden_activ_out_h001_004    tia_h_in_002_005-    120997.90407537823
Rh002_005_005+    hidden_activ_out_h001_005    tia_h_in_002_005+    119983.0173326794
Rh002_005_005-    hidden_activ_out_h001_005    tia_h_in_002_005-    120000
Rh002_006_005+    hidden_activ_out_h001_006    tia_h_in_002_005+    118649.9591637305
Rh002_006_005-    hidden_activ_out_h001_006    tia_h_in_002_005-    38865.46827086198
Rh002_007_005+    hidden_activ_out_h001_007    tia_h_in_002_005+    119542.23258003875
Rh002_007_005-    hidden_activ_out_h001_007    tia_h_in_002_005-    25712.178268768923
Rh002_008_005+    hidden_activ_out_h001_008    tia_h_in_002_005+    119195.72011416264
Rh002_008_005-    hidden_activ_out_h001_008    tia_h_in_002_005-    19801.478278833034
Rh002_009_005+    hidden_activ_out_h001_009    tia_h_in_002_005+    118854.10788789322
Rh002_009_005-    hidden_activ_out_h001_009    tia_h_in_002_005-    43972.05080098318
Rh002_010_005+    hidden_activ_out_h001_010    tia_h_in_002_005+    119621.48400469171
Rh002_010_005-    hidden_activ_out_h001_010    tia_h_in_002_005-    71008.09504950859
Rh002_011_005+    hidden_activ_out_h001_011    tia_h_in_002_005+    119531.97319784667
Rh002_011_005-    hidden_activ_out_h001_011    tia_h_in_002_005-    5000
Rh002_012_005+    hidden_activ_out_h001_012    tia_h_in_002_005+    120319.19927019638
Rh002_012_005-    hidden_activ_out_h001_012    tia_h_in_002_005-    76640.89029824715
Rh002_013_005+    hidden_activ_out_h001_013    tia_h_in_002_005+    118978.61146489413
Rh002_013_005-    hidden_activ_out_h001_013    tia_h_in_002_005-    29374.984558425167
Rh002_014_005+    hidden_activ_out_h001_014    tia_h_in_002_005+    91686.37564549557
Rh002_014_005-    hidden_activ_out_h001_014    tia_h_in_002_005-    121423.76774155513
Rh002_015_005+    hidden_activ_out_h001_015    tia_h_in_002_005+    121103.07715749885
Rh002_015_005-    hidden_activ_out_h001_015    tia_h_in_002_005-    47499.29266644817
Rh002_016_005+    hidden_activ_out_h001_016    tia_h_in_002_005+    16382.201894212027
Rh002_016_005-    hidden_activ_out_h001_016    tia_h_in_002_005-    121193.75601544506
Rh002_017_005+    hidden_activ_out_h001_017    tia_h_in_002_005+    26975.138652337107
Rh002_017_005-    hidden_activ_out_h001_017    tia_h_in_002_005-    119982.10313101015
Rh002_018_005+    hidden_activ_out_h001_018    tia_h_in_002_005+    119535.61228879365
Rh002_018_005-    hidden_activ_out_h001_018    tia_h_in_002_005-    66339.87927322071
Rh002_019_005+    hidden_activ_out_h001_019    tia_h_in_002_005+    120000
Rh002_019_005-    hidden_activ_out_h001_019    tia_h_in_002_005-    117779.8027773943
Rh002_020_005+    hidden_activ_out_h001_020    tia_h_in_002_005+    90673.34214787418
Rh002_020_005-    hidden_activ_out_h001_020    tia_h_in_002_005-    119897.0799702362

* Neuron 6
Rh002_001_006+    hidden_activ_out_h001_001    tia_h_in_002_006+    119806.97320802475
Rh002_001_006-    hidden_activ_out_h001_001    tia_h_in_002_006-    120000
Rh002_002_006+    hidden_activ_out_h001_002    tia_h_in_002_006+    41905.422646891355
Rh002_002_006-    hidden_activ_out_h001_002    tia_h_in_002_006-    120762.12027476955
Rh002_003_006+    hidden_activ_out_h001_003    tia_h_in_002_006+    121216.08713381732
Rh002_003_006-    hidden_activ_out_h001_003    tia_h_in_002_006-    5999.389881123192
Rh002_004_006+    hidden_activ_out_h001_004    tia_h_in_002_006+    119185.04910708636
Rh002_004_006-    hidden_activ_out_h001_004    tia_h_in_002_006-    102352.53583365296
Rh002_005_006+    hidden_activ_out_h001_005    tia_h_in_002_006+    6865.936414763047
Rh002_005_006-    hidden_activ_out_h001_005    tia_h_in_002_006-    120728.05258270237
Rh002_006_006+    hidden_activ_out_h001_006    tia_h_in_002_006+    100813.85156353071
Rh002_006_006-    hidden_activ_out_h001_006    tia_h_in_002_006-    120917.2830671943
Rh002_007_006+    hidden_activ_out_h001_007    tia_h_in_002_006+    25144.87795970538
Rh002_007_006-    hidden_activ_out_h001_007    tia_h_in_002_006-    120254.634626977
Rh002_008_006+    hidden_activ_out_h001_008    tia_h_in_002_006+    7879.48790760932
Rh002_008_006-    hidden_activ_out_h001_008    tia_h_in_002_006-    117746.31425816096
Rh002_009_006+    hidden_activ_out_h001_009    tia_h_in_002_006+    28632.75089961869
Rh002_009_006-    hidden_activ_out_h001_009    tia_h_in_002_006-    121357.23469085139
Rh002_010_006+    hidden_activ_out_h001_010    tia_h_in_002_006+    119355.5325258465
Rh002_010_006-    hidden_activ_out_h001_010    tia_h_in_002_006-    55504.45568494061
Rh002_011_006+    hidden_activ_out_h001_011    tia_h_in_002_006+    15121.689066448282
Rh002_011_006-    hidden_activ_out_h001_011    tia_h_in_002_006-    119163.47540920279
Rh002_012_006+    hidden_activ_out_h001_012    tia_h_in_002_006+    119360.8587752762
Rh002_012_006-    hidden_activ_out_h001_012    tia_h_in_002_006-    64487.59924051003
Rh002_013_006+    hidden_activ_out_h001_013    tia_h_in_002_006+    14845.761454117046
Rh002_013_006-    hidden_activ_out_h001_013    tia_h_in_002_006-    120434.13629192988
Rh002_014_006+    hidden_activ_out_h001_014    tia_h_in_002_006+    84506.07298792897
Rh002_014_006-    hidden_activ_out_h001_014    tia_h_in_002_006-    119169.31742526461
Rh002_015_006+    hidden_activ_out_h001_015    tia_h_in_002_006+    121040.17973047205
Rh002_015_006-    hidden_activ_out_h001_015    tia_h_in_002_006-    112678.45090071263
Rh002_016_006+    hidden_activ_out_h001_016    tia_h_in_002_006+    118529.18504126277
Rh002_016_006-    hidden_activ_out_h001_016    tia_h_in_002_006-    120000
Rh002_017_006+    hidden_activ_out_h001_017    tia_h_in_002_006+    5000
Rh002_017_006-    hidden_activ_out_h001_017    tia_h_in_002_006-    12550.464919424427
Rh002_018_006+    hidden_activ_out_h001_018    tia_h_in_002_006+    19129.34443266239
Rh002_018_006-    hidden_activ_out_h001_018    tia_h_in_002_006-    119392.91568925478
Rh002_019_006+    hidden_activ_out_h001_019    tia_h_in_002_006+    120792.23728693479
Rh002_019_006-    hidden_activ_out_h001_019    tia_h_in_002_006-    5165.972796755012
Rh002_020_006+    hidden_activ_out_h001_020    tia_h_in_002_006+    120379.2362364863
Rh002_020_006-    hidden_activ_out_h001_020    tia_h_in_002_006-    120000

* Neuron 7
Rh002_001_007+    hidden_activ_out_h001_001    tia_h_in_002_007+    28195.05700940881
Rh002_001_007-    hidden_activ_out_h001_001    tia_h_in_002_007-    120960.25957340485
Rh002_002_007+    hidden_activ_out_h001_002    tia_h_in_002_007+    120421.08011840843
Rh002_002_007-    hidden_activ_out_h001_002    tia_h_in_002_007-    9592.630065606721
Rh002_003_007+    hidden_activ_out_h001_003    tia_h_in_002_007+    120000
Rh002_003_007-    hidden_activ_out_h001_003    tia_h_in_002_007-    120676.4227595781
Rh002_004_007+    hidden_activ_out_h001_004    tia_h_in_002_007+    119487.6455338742
Rh002_004_007-    hidden_activ_out_h001_004    tia_h_in_002_007-    5000
Rh002_005_007+    hidden_activ_out_h001_005    tia_h_in_002_007+    118897.84075328174
Rh002_005_007-    hidden_activ_out_h001_005    tia_h_in_002_007-    120000
Rh002_006_007+    hidden_activ_out_h001_006    tia_h_in_002_007+    121547.14797310799
Rh002_006_007-    hidden_activ_out_h001_006    tia_h_in_002_007-    65338.68504501388
Rh002_007_007+    hidden_activ_out_h001_007    tia_h_in_002_007+    120187.01065381734
Rh002_007_007-    hidden_activ_out_h001_007    tia_h_in_002_007-    15096.600678487743
Rh002_008_007+    hidden_activ_out_h001_008    tia_h_in_002_007+    119670.56581579956
Rh002_008_007-    hidden_activ_out_h001_008    tia_h_in_002_007-    18748.282935013416
Rh002_009_007+    hidden_activ_out_h001_009    tia_h_in_002_007+    119106.81513344405
Rh002_009_007-    hidden_activ_out_h001_009    tia_h_in_002_007-    15266.835295813518
Rh002_010_007+    hidden_activ_out_h001_010    tia_h_in_002_007+    38693.65816154094
Rh002_010_007-    hidden_activ_out_h001_010    tia_h_in_002_007-    120259.20468180993
Rh002_011_007+    hidden_activ_out_h001_011    tia_h_in_002_007+    121791.00700957254
Rh002_011_007-    hidden_activ_out_h001_011    tia_h_in_002_007-    12139.536156814924
Rh002_012_007+    hidden_activ_out_h001_012    tia_h_in_002_007+    119128.42811689457
Rh002_012_007-    hidden_activ_out_h001_012    tia_h_in_002_007-    29615.721811309308
Rh002_013_007+    hidden_activ_out_h001_013    tia_h_in_002_007+    121002.96776731868
Rh002_013_007-    hidden_activ_out_h001_013    tia_h_in_002_007-    11035.380929369978
Rh002_014_007+    hidden_activ_out_h001_014    tia_h_in_002_007+    51126.23742664372
Rh002_014_007-    hidden_activ_out_h001_014    tia_h_in_002_007-    120775.00963181542
Rh002_015_007+    hidden_activ_out_h001_015    tia_h_in_002_007+    119512.10969736612
Rh002_015_007-    hidden_activ_out_h001_015    tia_h_in_002_007-    43250.35125933993
Rh002_016_007+    hidden_activ_out_h001_016    tia_h_in_002_007+    23237.43876624158
Rh002_016_007-    hidden_activ_out_h001_016    tia_h_in_002_007-    120000
Rh002_017_007+    hidden_activ_out_h001_017    tia_h_in_002_007+    85102.83373617113
Rh002_017_007-    hidden_activ_out_h001_017    tia_h_in_002_007-    120100.33524658947
Rh002_018_007+    hidden_activ_out_h001_018    tia_h_in_002_007+    121536.48243545838
Rh002_018_007-    hidden_activ_out_h001_018    tia_h_in_002_007-    25260.69331067818
Rh002_019_007+    hidden_activ_out_h001_019    tia_h_in_002_007+    20364.121626193228
Rh002_019_007-    hidden_activ_out_h001_019    tia_h_in_002_007-    121035.79686348712
Rh002_020_007+    hidden_activ_out_h001_020    tia_h_in_002_007+    120000
Rh002_020_007-    hidden_activ_out_h001_020    tia_h_in_002_007-    51773.959619134825

* Neuron 8
Rh002_001_008+    hidden_activ_out_h001_001    tia_h_in_002_008+    90023.43983624055
Rh002_001_008-    hidden_activ_out_h001_001    tia_h_in_002_008-    119481.36044874466
Rh002_002_008+    hidden_activ_out_h001_002    tia_h_in_002_008+    120568.52660164874
Rh002_002_008-    hidden_activ_out_h001_002    tia_h_in_002_008-    5656.617930582286
Rh002_003_008+    hidden_activ_out_h001_003    tia_h_in_002_008+    24145.873793320865
Rh002_003_008-    hidden_activ_out_h001_003    tia_h_in_002_008-    120151.62770159144
Rh002_004_008+    hidden_activ_out_h001_004    tia_h_in_002_008+    62702.34658024195
Rh002_004_008-    hidden_activ_out_h001_004    tia_h_in_002_008-    118923.29542081969
Rh002_005_008+    hidden_activ_out_h001_005    tia_h_in_002_008+    119418.97049043313
Rh002_005_008-    hidden_activ_out_h001_005    tia_h_in_002_008-    11809.898458325291
Rh002_006_008+    hidden_activ_out_h001_006    tia_h_in_002_008+    120361.32462459092
Rh002_006_008-    hidden_activ_out_h001_006    tia_h_in_002_008-    63375.15234944889
Rh002_007_008+    hidden_activ_out_h001_007    tia_h_in_002_008+    121223.74075948038
Rh002_007_008-    hidden_activ_out_h001_007    tia_h_in_002_008-    9254.237305982351
Rh002_008_008+    hidden_activ_out_h001_008    tia_h_in_002_008+    118481.61114425212
Rh002_008_008-    hidden_activ_out_h001_008    tia_h_in_002_008-    11848.590127195535
Rh002_009_008+    hidden_activ_out_h001_009    tia_h_in_002_008+    122444.88376563459
Rh002_009_008-    hidden_activ_out_h001_009    tia_h_in_002_008-    7099.803833780345
Rh002_010_008+    hidden_activ_out_h001_010    tia_h_in_002_008+    39190.02787917148
Rh002_010_008-    hidden_activ_out_h001_010    tia_h_in_002_008-    119842.67389110738
Rh002_011_008+    hidden_activ_out_h001_011    tia_h_in_002_008+    120567.13989250195
Rh002_011_008-    hidden_activ_out_h001_011    tia_h_in_002_008-    11523.886942742396
Rh002_012_008+    hidden_activ_out_h001_012    tia_h_in_002_008+    119938.7635030475
Rh002_012_008-    hidden_activ_out_h001_012    tia_h_in_002_008-    11551.405624383386
Rh002_013_008+    hidden_activ_out_h001_013    tia_h_in_002_008+    119536.82542060432
Rh002_013_008-    hidden_activ_out_h001_013    tia_h_in_002_008-    8561.569363843735
Rh002_014_008+    hidden_activ_out_h001_014    tia_h_in_002_008+    71657.20289858142
Rh002_014_008-    hidden_activ_out_h001_014    tia_h_in_002_008-    120671.56424445295
Rh002_015_008+    hidden_activ_out_h001_015    tia_h_in_002_008+    44606.20677169488
Rh002_015_008-    hidden_activ_out_h001_015    tia_h_in_002_008-    121194.2369299505
Rh002_016_008+    hidden_activ_out_h001_016    tia_h_in_002_008+    119973.95645158607
Rh002_016_008-    hidden_activ_out_h001_016    tia_h_in_002_008-    99784.71261407598
Rh002_017_008+    hidden_activ_out_h001_017    tia_h_in_002_008+    119852.31568194293
Rh002_017_008-    hidden_activ_out_h001_017    tia_h_in_002_008-    31099.428883429402
Rh002_018_008+    hidden_activ_out_h001_018    tia_h_in_002_008+    118825.57128231235
Rh002_018_008-    hidden_activ_out_h001_018    tia_h_in_002_008-    6451.550116160723
Rh002_019_008+    hidden_activ_out_h001_019    tia_h_in_002_008+    26050.582337465214
Rh002_019_008-    hidden_activ_out_h001_019    tia_h_in_002_008-    120000
Rh002_020_008+    hidden_activ_out_h001_020    tia_h_in_002_008+    120419.92312692085
Rh002_020_008-    hidden_activ_out_h001_020    tia_h_in_002_008-    7132.672126400319

* Neuron 9
Rh002_001_009+    hidden_activ_out_h001_001    tia_h_in_002_009+    109881.69925989857
Rh002_001_009-    hidden_activ_out_h001_001    tia_h_in_002_009-    119835.09196229295
Rh002_002_009+    hidden_activ_out_h001_002    tia_h_in_002_009+    120207.27647881092
Rh002_002_009-    hidden_activ_out_h001_002    tia_h_in_002_009-    8337.978263263058
Rh002_003_009+    hidden_activ_out_h001_003    tia_h_in_002_009+    16885.658713585493
Rh002_003_009-    hidden_activ_out_h001_003    tia_h_in_002_009-    121527.52044143678
Rh002_004_009+    hidden_activ_out_h001_004    tia_h_in_002_009+    120406.84606701524
Rh002_004_009-    hidden_activ_out_h001_004    tia_h_in_002_009-    82870.62469840697
Rh002_005_009+    hidden_activ_out_h001_005    tia_h_in_002_009+    119926.62995591245
Rh002_005_009-    hidden_activ_out_h001_005    tia_h_in_002_009-    9833.800811846544
Rh002_006_009+    hidden_activ_out_h001_006    tia_h_in_002_009+    41330.970737683034
Rh002_006_009-    hidden_activ_out_h001_006    tia_h_in_002_009-    119941.3333661719
Rh002_007_009+    hidden_activ_out_h001_007    tia_h_in_002_009+    119640.03455611206
Rh002_007_009-    hidden_activ_out_h001_007    tia_h_in_002_009-    12068.81207574109
Rh002_008_009+    hidden_activ_out_h001_008    tia_h_in_002_009+    5000
Rh002_008_009-    hidden_activ_out_h001_008    tia_h_in_002_009-    12591.959921504254
Rh002_009_009+    hidden_activ_out_h001_009    tia_h_in_002_009+    120437.83797291583
Rh002_009_009-    hidden_activ_out_h001_009    tia_h_in_002_009-    8875.137662122781
Rh002_010_009+    hidden_activ_out_h001_010    tia_h_in_002_009+    47681.06402041604
Rh002_010_009-    hidden_activ_out_h001_010    tia_h_in_002_009-    120408.06536501106
Rh002_011_009+    hidden_activ_out_h001_011    tia_h_in_002_009+    120000
Rh002_011_009-    hidden_activ_out_h001_011    tia_h_in_002_009-    10742.963911483102
Rh002_012_009+    hidden_activ_out_h001_012    tia_h_in_002_009+    5000
Rh002_012_009-    hidden_activ_out_h001_012    tia_h_in_002_009-    5000
Rh002_013_009+    hidden_activ_out_h001_013    tia_h_in_002_009+    120702.00556409956
Rh002_013_009-    hidden_activ_out_h001_013    tia_h_in_002_009-    7936.497126436874
Rh002_014_009+    hidden_activ_out_h001_014    tia_h_in_002_009+    62817.937216397244
Rh002_014_009-    hidden_activ_out_h001_014    tia_h_in_002_009-    120441.72548717697
Rh002_015_009+    hidden_activ_out_h001_015    tia_h_in_002_009+    120654.72838849983
Rh002_015_009-    hidden_activ_out_h001_015    tia_h_in_002_009-    110322.76606291205
Rh002_016_009+    hidden_activ_out_h001_016    tia_h_in_002_009+    121424.89544242629
Rh002_016_009-    hidden_activ_out_h001_016    tia_h_in_002_009-    120000
Rh002_017_009+    hidden_activ_out_h001_017    tia_h_in_002_009+    120652.38417709268
Rh002_017_009-    hidden_activ_out_h001_017    tia_h_in_002_009-    93080.4644318832
Rh002_018_009+    hidden_activ_out_h001_018    tia_h_in_002_009+    118494.57623689783
Rh002_018_009-    hidden_activ_out_h001_018    tia_h_in_002_009-    13358.289707301024
Rh002_019_009+    hidden_activ_out_h001_019    tia_h_in_002_009+    24903.776593336064
Rh002_019_009-    hidden_activ_out_h001_019    tia_h_in_002_009-    120115.59349285265
Rh002_020_009+    hidden_activ_out_h001_020    tia_h_in_002_009+    119427.06615231307
Rh002_020_009-    hidden_activ_out_h001_020    tia_h_in_002_009-    29558.534409320066

* Neuron 10
Rh002_001_010+    hidden_activ_out_h001_001    tia_h_in_002_010+    14082.899926172258
Rh002_001_010-    hidden_activ_out_h001_001    tia_h_in_002_010-    119086.06433855653
Rh002_002_010+    hidden_activ_out_h001_002    tia_h_in_002_010+    119370.7221083249
Rh002_002_010-    hidden_activ_out_h001_002    tia_h_in_002_010-    5000
Rh002_003_010+    hidden_activ_out_h001_003    tia_h_in_002_010+    19609.57348282995
Rh002_003_010-    hidden_activ_out_h001_003    tia_h_in_002_010-    120526.25791375857
Rh002_004_010+    hidden_activ_out_h001_004    tia_h_in_002_010+    49470.27955701535
Rh002_004_010-    hidden_activ_out_h001_004    tia_h_in_002_010-    5000
Rh002_005_010+    hidden_activ_out_h001_005    tia_h_in_002_010+    119563.81037027939
Rh002_005_010-    hidden_activ_out_h001_005    tia_h_in_002_010-    14610.232766612135
Rh002_006_010+    hidden_activ_out_h001_006    tia_h_in_002_010+    39750.96239240636
Rh002_006_010-    hidden_activ_out_h001_006    tia_h_in_002_010-    121009.41460840001
Rh002_007_010+    hidden_activ_out_h001_007    tia_h_in_002_010+    119961.88300216745
Rh002_007_010-    hidden_activ_out_h001_007    tia_h_in_002_010-    24493.79230780017
Rh002_008_010+    hidden_activ_out_h001_008    tia_h_in_002_010+    119401.38055323425
Rh002_008_010-    hidden_activ_out_h001_008    tia_h_in_002_010-    17750.27413027818
Rh002_009_010+    hidden_activ_out_h001_009    tia_h_in_002_010+    120963.91941707788
Rh002_009_010-    hidden_activ_out_h001_009    tia_h_in_002_010-    40144.881998347904
Rh002_010_010+    hidden_activ_out_h001_010    tia_h_in_002_010+    120172.57231899195
Rh002_010_010-    hidden_activ_out_h001_010    tia_h_in_002_010-    48402.56778440959
Rh002_011_010+    hidden_activ_out_h001_011    tia_h_in_002_010+    120531.24893394703
Rh002_011_010-    hidden_activ_out_h001_011    tia_h_in_002_010-    24980.80499811087
Rh002_012_010+    hidden_activ_out_h001_012    tia_h_in_002_010+    119678.11082344284
Rh002_012_010-    hidden_activ_out_h001_012    tia_h_in_002_010-    71293.81012976891
Rh002_013_010+    hidden_activ_out_h001_013    tia_h_in_002_010+    119327.46140238376
Rh002_013_010-    hidden_activ_out_h001_013    tia_h_in_002_010-    30510.11636458869
Rh002_014_010+    hidden_activ_out_h001_014    tia_h_in_002_010+    97071.74208091269
Rh002_014_010-    hidden_activ_out_h001_014    tia_h_in_002_010-    5000
Rh002_015_010+    hidden_activ_out_h001_015    tia_h_in_002_010+    52403.86059571801
Rh002_015_010-    hidden_activ_out_h001_015    tia_h_in_002_010-    119413.35865730407
Rh002_016_010+    hidden_activ_out_h001_016    tia_h_in_002_010+    13940.147828464455
Rh002_016_010-    hidden_activ_out_h001_016    tia_h_in_002_010-    122518.15321274151
Rh002_017_010+    hidden_activ_out_h001_017    tia_h_in_002_010+    22300.79600653302
Rh002_017_010-    hidden_activ_out_h001_017    tia_h_in_002_010-    118210.88796601082
Rh002_018_010+    hidden_activ_out_h001_018    tia_h_in_002_010+    120029.24625528046
Rh002_018_010-    hidden_activ_out_h001_018    tia_h_in_002_010-    66045.27280834335
Rh002_019_010+    hidden_activ_out_h001_019    tia_h_in_002_010+    5000
Rh002_019_010-    hidden_activ_out_h001_019    tia_h_in_002_010-    5000
Rh002_020_010+    hidden_activ_out_h001_020    tia_h_in_002_010+    106218.67069807915
Rh002_020_010-    hidden_activ_out_h001_020    tia_h_in_002_010-    5000

* ----- Bias
    
        
Rb_h002_001+    b_002    tia_h_in_002_001+    42564.60949032792
Rb_h002_001-    b_002    tia_h_in_002_001-    120392.21536573823
Rb_h002_002+    b_002    tia_h_in_002_002+    33420.586003557575
Rb_h002_002-    b_002    tia_h_in_002_002-    120733.07795649106
Rb_h002_003+    b_002    tia_h_in_002_003+    31079.36694168635
Rb_h002_003-    b_002    tia_h_in_002_003-    120178.32283734417
Rb_h002_004+    b_002    tia_h_in_002_004+    61985.248106708954
Rb_h002_004-    b_002    tia_h_in_002_004-    119018.96106908204
Rb_h002_005+    b_002    tia_h_in_002_005+    60993.71925548039
Rb_h002_005-    b_002    tia_h_in_002_005-    120194.16281542076
Rb_h002_006+    b_002    tia_h_in_002_006+    43666.877571620855
Rb_h002_006-    b_002    tia_h_in_002_006-    120267.53272148679
Rb_h002_007+    b_002    tia_h_in_002_007+    32074.149354544003
Rb_h002_007-    b_002    tia_h_in_002_007-    119726.04714714253
Rb_h002_008+    b_002    tia_h_in_002_008+    25889.898074505887
Rb_h002_008-    b_002    tia_h_in_002_008-    121178.58002246462
Rb_h002_009+    b_002    tia_h_in_002_009+    27926.727171194678
Rb_h002_009-    b_002    tia_h_in_002_009-    119307.70487537142
Rb_h002_010+    b_002    tia_h_in_002_010+    59253.044724839485
Rb_h002_010-    b_002    tia_h_in_002_010-    120729.4665676119

* ----- Weights
* Layer 003

* Neuron 1
Rh003_001_001+    hidden_activ_out_h002_001    tia_h_in_003_001+    5000
Rh003_001_001-    hidden_activ_out_h002_001    tia_h_in_003_001-    5961.259916061574
Rh003_002_001+    hidden_activ_out_h002_002    tia_h_in_003_001+    4983.723487476977
Rh003_002_001-    hidden_activ_out_h002_002    tia_h_in_003_001-    120252.21884275884
Rh003_003_001+    hidden_activ_out_h002_003    tia_h_in_003_001+    120000
Rh003_003_001-    hidden_activ_out_h002_003    tia_h_in_003_001-    118403.92900070558
Rh003_004_001+    hidden_activ_out_h002_004    tia_h_in_003_001+    14143.80523067764
Rh003_004_001-    hidden_activ_out_h002_004    tia_h_in_003_001-    120000
Rh003_005_001+    hidden_activ_out_h002_005    tia_h_in_003_001+    11149.708350336226
Rh003_005_001-    hidden_activ_out_h002_005    tia_h_in_003_001-    121246.0720726309
Rh003_006_001+    hidden_activ_out_h002_006    tia_h_in_003_001+    119563.6888382225
Rh003_006_001-    hidden_activ_out_h002_006    tia_h_in_003_001-    5781.782644360064
Rh003_007_001+    hidden_activ_out_h002_007    tia_h_in_003_001+    9266.84158933853
Rh003_007_001-    hidden_activ_out_h002_007    tia_h_in_003_001-    118231.19582345875
Rh003_008_001+    hidden_activ_out_h002_008    tia_h_in_003_001+    6089.438317136861
Rh003_008_001-    hidden_activ_out_h002_008    tia_h_in_003_001-    120029.13036135715
Rh003_009_001+    hidden_activ_out_h002_009    tia_h_in_003_001+    7204.182871594563
Rh003_009_001-    hidden_activ_out_h002_009    tia_h_in_003_001-    120276.36107510292
Rh003_010_001+    hidden_activ_out_h002_010    tia_h_in_003_001+    12638.392244634002
Rh003_010_001-    hidden_activ_out_h002_010    tia_h_in_003_001-    120093.09666317259

* ----- Bias
    
        
Rb_h003_001+    b_003    tia_h_in_003_001+    118512.32188555584
Rb_h003_001-    b_003    tia_h_in_003_001-    7641.237111119246


* ----- Difference (V(R+) - V(R-))

* Layer 000
* Neuron 1
Rh001_fb_001+     tia_h_in_001_001+ tia_h_out_001_001+ 4785.331062648607
Rh001_fb_001-     tia_h_in_001_001- tia_h_out_001_001- 4785.331062648607
XUh001_001+       0 tia_h_in_001_001+ Vcc+ Vcc- tia_h_out_001_001+ Ve OPA684_0
XUh001_001-       0 tia_h_in_001_001- Vcc+ Vcc- tia_h_out_001_001- Ve OPA684_0
Rh001_sum_001+    tia_h_out_001_001+ sum_h_in_001_001- 260
Rh001_sum_001-    tia_h_out_001_001- sum_h_in_001_001+ 260
Rh001_sum_l_001   sum_h_in_001_001+ 0 650.0
Rh001_sum_fb_001  sum_h_in_001_001- sum_h_out_001_001 650.0
XUh001_sum_001    sum_h_in_001_001+ sum_h_in_001_001- Vcc+ Vcc- sum_h_out_001_001 MAX4223
* Neuron 2
Rh001_fb_002+     tia_h_in_001_002+ tia_h_out_001_002+ 4785.331062648607
Rh001_fb_002-     tia_h_in_001_002- tia_h_out_001_002- 4785.331062648607
XUh001_002+       0 tia_h_in_001_002+ Vcc+ Vcc- tia_h_out_001_002+ Ve OPA684_0
XUh001_002-       0 tia_h_in_001_002- Vcc+ Vcc- tia_h_out_001_002- Ve OPA684_0
Rh001_sum_002+    tia_h_out_001_002+ sum_h_in_001_002- 260
Rh001_sum_002-    tia_h_out_001_002- sum_h_in_001_002+ 260
Rh001_sum_l_002   sum_h_in_001_002+ 0 650.0
Rh001_sum_fb_002  sum_h_in_001_002- sum_h_out_001_002 650.0
XUh001_sum_002    sum_h_in_001_002+ sum_h_in_001_002- Vcc+ Vcc- sum_h_out_001_002 MAX4223
* Neuron 3
Rh001_fb_003+     tia_h_in_001_003+ tia_h_out_001_003+ 4785.331062648607
Rh001_fb_003-     tia_h_in_001_003- tia_h_out_001_003- 4785.331062648607
XUh001_003+       0 tia_h_in_001_003+ Vcc+ Vcc- tia_h_out_001_003+ Ve OPA684_0
XUh001_003-       0 tia_h_in_001_003- Vcc+ Vcc- tia_h_out_001_003- Ve OPA684_0
Rh001_sum_003+    tia_h_out_001_003+ sum_h_in_001_003- 260
Rh001_sum_003-    tia_h_out_001_003- sum_h_in_001_003+ 260
Rh001_sum_l_003   sum_h_in_001_003+ 0 650.0
Rh001_sum_fb_003  sum_h_in_001_003- sum_h_out_001_003 650.0
XUh001_sum_003    sum_h_in_001_003+ sum_h_in_001_003- Vcc+ Vcc- sum_h_out_001_003 MAX4223
* Neuron 4
Rh001_fb_004+     tia_h_in_001_004+ tia_h_out_001_004+ 4785.331062648607
Rh001_fb_004-     tia_h_in_001_004- tia_h_out_001_004- 4785.331062648607
XUh001_004+       0 tia_h_in_001_004+ Vcc+ Vcc- tia_h_out_001_004+ Ve OPA684_0
XUh001_004-       0 tia_h_in_001_004- Vcc+ Vcc- tia_h_out_001_004- Ve OPA684_0
Rh001_sum_004+    tia_h_out_001_004+ sum_h_in_001_004- 260
Rh001_sum_004-    tia_h_out_001_004- sum_h_in_001_004+ 260
Rh001_sum_l_004   sum_h_in_001_004+ 0 650.0
Rh001_sum_fb_004  sum_h_in_001_004- sum_h_out_001_004 650.0
XUh001_sum_004    sum_h_in_001_004+ sum_h_in_001_004- Vcc+ Vcc- sum_h_out_001_004 MAX4223
* Neuron 5
Rh001_fb_005+     tia_h_in_001_005+ tia_h_out_001_005+ 4785.331062648607
Rh001_fb_005-     tia_h_in_001_005- tia_h_out_001_005- 4785.331062648607
XUh001_005+       0 tia_h_in_001_005+ Vcc+ Vcc- tia_h_out_001_005+ Ve OPA684_0
XUh001_005-       0 tia_h_in_001_005- Vcc+ Vcc- tia_h_out_001_005- Ve OPA684_0
Rh001_sum_005+    tia_h_out_001_005+ sum_h_in_001_005- 260
Rh001_sum_005-    tia_h_out_001_005- sum_h_in_001_005+ 260
Rh001_sum_l_005   sum_h_in_001_005+ 0 650.0
Rh001_sum_fb_005  sum_h_in_001_005- sum_h_out_001_005 650.0
XUh001_sum_005    sum_h_in_001_005+ sum_h_in_001_005- Vcc+ Vcc- sum_h_out_001_005 MAX4223
* Neuron 6
Rh001_fb_006+     tia_h_in_001_006+ tia_h_out_001_006+ 4785.331062648607
Rh001_fb_006-     tia_h_in_001_006- tia_h_out_001_006- 4785.331062648607
XUh001_006+       0 tia_h_in_001_006+ Vcc+ Vcc- tia_h_out_001_006+ Ve OPA684_0
XUh001_006-       0 tia_h_in_001_006- Vcc+ Vcc- tia_h_out_001_006- Ve OPA684_0
Rh001_sum_006+    tia_h_out_001_006+ sum_h_in_001_006- 260
Rh001_sum_006-    tia_h_out_001_006- sum_h_in_001_006+ 260
Rh001_sum_l_006   sum_h_in_001_006+ 0 650.0
Rh001_sum_fb_006  sum_h_in_001_006- sum_h_out_001_006 650.0
XUh001_sum_006    sum_h_in_001_006+ sum_h_in_001_006- Vcc+ Vcc- sum_h_out_001_006 MAX4223
* Neuron 7
Rh001_fb_007+     tia_h_in_001_007+ tia_h_out_001_007+ 4785.331062648607
Rh001_fb_007-     tia_h_in_001_007- tia_h_out_001_007- 4785.331062648607
XUh001_007+       0 tia_h_in_001_007+ Vcc+ Vcc- tia_h_out_001_007+ Ve OPA684_0
XUh001_007-       0 tia_h_in_001_007- Vcc+ Vcc- tia_h_out_001_007- Ve OPA684_0
Rh001_sum_007+    tia_h_out_001_007+ sum_h_in_001_007- 260
Rh001_sum_007-    tia_h_out_001_007- sum_h_in_001_007+ 260
Rh001_sum_l_007   sum_h_in_001_007+ 0 650.0
Rh001_sum_fb_007  sum_h_in_001_007- sum_h_out_001_007 650.0
XUh001_sum_007    sum_h_in_001_007+ sum_h_in_001_007- Vcc+ Vcc- sum_h_out_001_007 MAX4223
* Neuron 8
Rh001_fb_008+     tia_h_in_001_008+ tia_h_out_001_008+ 4785.331062648607
Rh001_fb_008-     tia_h_in_001_008- tia_h_out_001_008- 4785.331062648607
XUh001_008+       0 tia_h_in_001_008+ Vcc+ Vcc- tia_h_out_001_008+ Ve OPA684_0
XUh001_008-       0 tia_h_in_001_008- Vcc+ Vcc- tia_h_out_001_008- Ve OPA684_0
Rh001_sum_008+    tia_h_out_001_008+ sum_h_in_001_008- 260
Rh001_sum_008-    tia_h_out_001_008- sum_h_in_001_008+ 260
Rh001_sum_l_008   sum_h_in_001_008+ 0 650.0
Rh001_sum_fb_008  sum_h_in_001_008- sum_h_out_001_008 650.0
XUh001_sum_008    sum_h_in_001_008+ sum_h_in_001_008- Vcc+ Vcc- sum_h_out_001_008 MAX4223
* Neuron 9
Rh001_fb_009+     tia_h_in_001_009+ tia_h_out_001_009+ 4785.331062648607
Rh001_fb_009-     tia_h_in_001_009- tia_h_out_001_009- 4785.331062648607
XUh001_009+       0 tia_h_in_001_009+ Vcc+ Vcc- tia_h_out_001_009+ Ve OPA684_0
XUh001_009-       0 tia_h_in_001_009- Vcc+ Vcc- tia_h_out_001_009- Ve OPA684_0
Rh001_sum_009+    tia_h_out_001_009+ sum_h_in_001_009- 260
Rh001_sum_009-    tia_h_out_001_009- sum_h_in_001_009+ 260
Rh001_sum_l_009   sum_h_in_001_009+ 0 650.0
Rh001_sum_fb_009  sum_h_in_001_009- sum_h_out_001_009 650.0
XUh001_sum_009    sum_h_in_001_009+ sum_h_in_001_009- Vcc+ Vcc- sum_h_out_001_009 MAX4223
* Neuron 10
Rh001_fb_010+     tia_h_in_001_010+ tia_h_out_001_010+ 4785.331062648607
Rh001_fb_010-     tia_h_in_001_010- tia_h_out_001_010- 4785.331062648607
XUh001_010+       0 tia_h_in_001_010+ Vcc+ Vcc- tia_h_out_001_010+ Ve OPA684_0
XUh001_010-       0 tia_h_in_001_010- Vcc+ Vcc- tia_h_out_001_010- Ve OPA684_0
Rh001_sum_010+    tia_h_out_001_010+ sum_h_in_001_010- 260
Rh001_sum_010-    tia_h_out_001_010- sum_h_in_001_010+ 260
Rh001_sum_l_010   sum_h_in_001_010+ 0 650.0
Rh001_sum_fb_010  sum_h_in_001_010- sum_h_out_001_010 650.0
XUh001_sum_010    sum_h_in_001_010+ sum_h_in_001_010- Vcc+ Vcc- sum_h_out_001_010 MAX4223
* Neuron 11
Rh001_fb_011+     tia_h_in_001_011+ tia_h_out_001_011+ 4785.331062648607
Rh001_fb_011-     tia_h_in_001_011- tia_h_out_001_011- 4785.331062648607
XUh001_011+       0 tia_h_in_001_011+ Vcc+ Vcc- tia_h_out_001_011+ Ve OPA684_0
XUh001_011-       0 tia_h_in_001_011- Vcc+ Vcc- tia_h_out_001_011- Ve OPA684_0
Rh001_sum_011+    tia_h_out_001_011+ sum_h_in_001_011- 260
Rh001_sum_011-    tia_h_out_001_011- sum_h_in_001_011+ 260
Rh001_sum_l_011   sum_h_in_001_011+ 0 650.0
Rh001_sum_fb_011  sum_h_in_001_011- sum_h_out_001_011 650.0
XUh001_sum_011    sum_h_in_001_011+ sum_h_in_001_011- Vcc+ Vcc- sum_h_out_001_011 MAX4223
* Neuron 12
Rh001_fb_012+     tia_h_in_001_012+ tia_h_out_001_012+ 4785.331062648607
Rh001_fb_012-     tia_h_in_001_012- tia_h_out_001_012- 4785.331062648607
XUh001_012+       0 tia_h_in_001_012+ Vcc+ Vcc- tia_h_out_001_012+ Ve OPA684_0
XUh001_012-       0 tia_h_in_001_012- Vcc+ Vcc- tia_h_out_001_012- Ve OPA684_0
Rh001_sum_012+    tia_h_out_001_012+ sum_h_in_001_012- 260
Rh001_sum_012-    tia_h_out_001_012- sum_h_in_001_012+ 260
Rh001_sum_l_012   sum_h_in_001_012+ 0 650.0
Rh001_sum_fb_012  sum_h_in_001_012- sum_h_out_001_012 650.0
XUh001_sum_012    sum_h_in_001_012+ sum_h_in_001_012- Vcc+ Vcc- sum_h_out_001_012 MAX4223
* Neuron 13
Rh001_fb_013+     tia_h_in_001_013+ tia_h_out_001_013+ 4785.331062648607
Rh001_fb_013-     tia_h_in_001_013- tia_h_out_001_013- 4785.331062648607
XUh001_013+       0 tia_h_in_001_013+ Vcc+ Vcc- tia_h_out_001_013+ Ve OPA684_0
XUh001_013-       0 tia_h_in_001_013- Vcc+ Vcc- tia_h_out_001_013- Ve OPA684_0
Rh001_sum_013+    tia_h_out_001_013+ sum_h_in_001_013- 260
Rh001_sum_013-    tia_h_out_001_013- sum_h_in_001_013+ 260
Rh001_sum_l_013   sum_h_in_001_013+ 0 650.0
Rh001_sum_fb_013  sum_h_in_001_013- sum_h_out_001_013 650.0
XUh001_sum_013    sum_h_in_001_013+ sum_h_in_001_013- Vcc+ Vcc- sum_h_out_001_013 MAX4223
* Neuron 14
Rh001_fb_014+     tia_h_in_001_014+ tia_h_out_001_014+ 4785.331062648607
Rh001_fb_014-     tia_h_in_001_014- tia_h_out_001_014- 4785.331062648607
XUh001_014+       0 tia_h_in_001_014+ Vcc+ Vcc- tia_h_out_001_014+ Ve OPA684_0
XUh001_014-       0 tia_h_in_001_014- Vcc+ Vcc- tia_h_out_001_014- Ve OPA684_0
Rh001_sum_014+    tia_h_out_001_014+ sum_h_in_001_014- 260
Rh001_sum_014-    tia_h_out_001_014- sum_h_in_001_014+ 260
Rh001_sum_l_014   sum_h_in_001_014+ 0 650.0
Rh001_sum_fb_014  sum_h_in_001_014- sum_h_out_001_014 650.0
XUh001_sum_014    sum_h_in_001_014+ sum_h_in_001_014- Vcc+ Vcc- sum_h_out_001_014 MAX4223
* Neuron 15
Rh001_fb_015+     tia_h_in_001_015+ tia_h_out_001_015+ 4785.331062648607
Rh001_fb_015-     tia_h_in_001_015- tia_h_out_001_015- 4785.331062648607
XUh001_015+       0 tia_h_in_001_015+ Vcc+ Vcc- tia_h_out_001_015+ Ve OPA684_0
XUh001_015-       0 tia_h_in_001_015- Vcc+ Vcc- tia_h_out_001_015- Ve OPA684_0
Rh001_sum_015+    tia_h_out_001_015+ sum_h_in_001_015- 260
Rh001_sum_015-    tia_h_out_001_015- sum_h_in_001_015+ 260
Rh001_sum_l_015   sum_h_in_001_015+ 0 650.0
Rh001_sum_fb_015  sum_h_in_001_015- sum_h_out_001_015 650.0
XUh001_sum_015    sum_h_in_001_015+ sum_h_in_001_015- Vcc+ Vcc- sum_h_out_001_015 MAX4223
* Neuron 16
Rh001_fb_016+     tia_h_in_001_016+ tia_h_out_001_016+ 4785.331062648607
Rh001_fb_016-     tia_h_in_001_016- tia_h_out_001_016- 4785.331062648607
XUh001_016+       0 tia_h_in_001_016+ Vcc+ Vcc- tia_h_out_001_016+ Ve OPA684_0
XUh001_016-       0 tia_h_in_001_016- Vcc+ Vcc- tia_h_out_001_016- Ve OPA684_0
Rh001_sum_016+    tia_h_out_001_016+ sum_h_in_001_016- 260
Rh001_sum_016-    tia_h_out_001_016- sum_h_in_001_016+ 260
Rh001_sum_l_016   sum_h_in_001_016+ 0 650.0
Rh001_sum_fb_016  sum_h_in_001_016- sum_h_out_001_016 650.0
XUh001_sum_016    sum_h_in_001_016+ sum_h_in_001_016- Vcc+ Vcc- sum_h_out_001_016 MAX4223
* Neuron 17
Rh001_fb_017+     tia_h_in_001_017+ tia_h_out_001_017+ 4785.331062648607
Rh001_fb_017-     tia_h_in_001_017- tia_h_out_001_017- 4785.331062648607
XUh001_017+       0 tia_h_in_001_017+ Vcc+ Vcc- tia_h_out_001_017+ Ve OPA684_0
XUh001_017-       0 tia_h_in_001_017- Vcc+ Vcc- tia_h_out_001_017- Ve OPA684_0
Rh001_sum_017+    tia_h_out_001_017+ sum_h_in_001_017- 260
Rh001_sum_017-    tia_h_out_001_017- sum_h_in_001_017+ 260
Rh001_sum_l_017   sum_h_in_001_017+ 0 650.0
Rh001_sum_fb_017  sum_h_in_001_017- sum_h_out_001_017 650.0
XUh001_sum_017    sum_h_in_001_017+ sum_h_in_001_017- Vcc+ Vcc- sum_h_out_001_017 MAX4223
* Neuron 18
Rh001_fb_018+     tia_h_in_001_018+ tia_h_out_001_018+ 4785.331062648607
Rh001_fb_018-     tia_h_in_001_018- tia_h_out_001_018- 4785.331062648607
XUh001_018+       0 tia_h_in_001_018+ Vcc+ Vcc- tia_h_out_001_018+ Ve OPA684_0
XUh001_018-       0 tia_h_in_001_018- Vcc+ Vcc- tia_h_out_001_018- Ve OPA684_0
Rh001_sum_018+    tia_h_out_001_018+ sum_h_in_001_018- 260
Rh001_sum_018-    tia_h_out_001_018- sum_h_in_001_018+ 260
Rh001_sum_l_018   sum_h_in_001_018+ 0 650.0
Rh001_sum_fb_018  sum_h_in_001_018- sum_h_out_001_018 650.0
XUh001_sum_018    sum_h_in_001_018+ sum_h_in_001_018- Vcc+ Vcc- sum_h_out_001_018 MAX4223
* Neuron 19
Rh001_fb_019+     tia_h_in_001_019+ tia_h_out_001_019+ 4785.331062648607
Rh001_fb_019-     tia_h_in_001_019- tia_h_out_001_019- 4785.331062648607
XUh001_019+       0 tia_h_in_001_019+ Vcc+ Vcc- tia_h_out_001_019+ Ve OPA684_0
XUh001_019-       0 tia_h_in_001_019- Vcc+ Vcc- tia_h_out_001_019- Ve OPA684_0
Rh001_sum_019+    tia_h_out_001_019+ sum_h_in_001_019- 260
Rh001_sum_019-    tia_h_out_001_019- sum_h_in_001_019+ 260
Rh001_sum_l_019   sum_h_in_001_019+ 0 650.0
Rh001_sum_fb_019  sum_h_in_001_019- sum_h_out_001_019 650.0
XUh001_sum_019    sum_h_in_001_019+ sum_h_in_001_019- Vcc+ Vcc- sum_h_out_001_019 MAX4223
* Neuron 20
Rh001_fb_020+     tia_h_in_001_020+ tia_h_out_001_020+ 4785.331062648607
Rh001_fb_020-     tia_h_in_001_020- tia_h_out_001_020- 4785.331062648607
XUh001_020+       0 tia_h_in_001_020+ Vcc+ Vcc- tia_h_out_001_020+ Ve OPA684_0
XUh001_020-       0 tia_h_in_001_020- Vcc+ Vcc- tia_h_out_001_020- Ve OPA684_0
Rh001_sum_020+    tia_h_out_001_020+ sum_h_in_001_020- 260
Rh001_sum_020-    tia_h_out_001_020- sum_h_in_001_020+ 260
Rh001_sum_l_020   sum_h_in_001_020+ 0 650.0
Rh001_sum_fb_020  sum_h_in_001_020- sum_h_out_001_020 650.0
XUh001_sum_020    sum_h_in_001_020+ sum_h_in_001_020- Vcc+ Vcc- sum_h_out_001_020 MAX4223

* Layer 001
* Neuron 1
Rh002_fb_001+     tia_h_in_002_001+ tia_h_out_002_001+ 4785.331062648607
Rh002_fb_001-     tia_h_in_002_001- tia_h_out_002_001- 4785.331062648607
XUh002_001+       0 tia_h_in_002_001+ Vcc+ Vcc- tia_h_out_002_001+ Ve OPA684_0
XUh002_001-       0 tia_h_in_002_001- Vcc+ Vcc- tia_h_out_002_001- Ve OPA684_0
Rh002_sum_001+    tia_h_out_002_001+ sum_h_in_002_001- 260
Rh002_sum_001-    tia_h_out_002_001- sum_h_in_002_001+ 260
Rh002_sum_l_001   sum_h_in_002_001+ 0 650.0
Rh002_sum_fb_001  sum_h_in_002_001- sum_h_out_002_001 650.0
XUh002_sum_001    sum_h_in_002_001+ sum_h_in_002_001- Vcc+ Vcc- sum_h_out_002_001 MAX4223
* Neuron 2
Rh002_fb_002+     tia_h_in_002_002+ tia_h_out_002_002+ 4785.331062648607
Rh002_fb_002-     tia_h_in_002_002- tia_h_out_002_002- 4785.331062648607
XUh002_002+       0 tia_h_in_002_002+ Vcc+ Vcc- tia_h_out_002_002+ Ve OPA684_0
XUh002_002-       0 tia_h_in_002_002- Vcc+ Vcc- tia_h_out_002_002- Ve OPA684_0
Rh002_sum_002+    tia_h_out_002_002+ sum_h_in_002_002- 260
Rh002_sum_002-    tia_h_out_002_002- sum_h_in_002_002+ 260
Rh002_sum_l_002   sum_h_in_002_002+ 0 650.0
Rh002_sum_fb_002  sum_h_in_002_002- sum_h_out_002_002 650.0
XUh002_sum_002    sum_h_in_002_002+ sum_h_in_002_002- Vcc+ Vcc- sum_h_out_002_002 MAX4223
* Neuron 3
Rh002_fb_003+     tia_h_in_002_003+ tia_h_out_002_003+ 4785.331062648607
Rh002_fb_003-     tia_h_in_002_003- tia_h_out_002_003- 4785.331062648607
XUh002_003+       0 tia_h_in_002_003+ Vcc+ Vcc- tia_h_out_002_003+ Ve OPA684_0
XUh002_003-       0 tia_h_in_002_003- Vcc+ Vcc- tia_h_out_002_003- Ve OPA684_0
Rh002_sum_003+    tia_h_out_002_003+ sum_h_in_002_003- 260
Rh002_sum_003-    tia_h_out_002_003- sum_h_in_002_003+ 260
Rh002_sum_l_003   sum_h_in_002_003+ 0 650.0
Rh002_sum_fb_003  sum_h_in_002_003- sum_h_out_002_003 650.0
XUh002_sum_003    sum_h_in_002_003+ sum_h_in_002_003- Vcc+ Vcc- sum_h_out_002_003 MAX4223
* Neuron 4
Rh002_fb_004+     tia_h_in_002_004+ tia_h_out_002_004+ 4785.331062648607
Rh002_fb_004-     tia_h_in_002_004- tia_h_out_002_004- 4785.331062648607
XUh002_004+       0 tia_h_in_002_004+ Vcc+ Vcc- tia_h_out_002_004+ Ve OPA684_0
XUh002_004-       0 tia_h_in_002_004- Vcc+ Vcc- tia_h_out_002_004- Ve OPA684_0
Rh002_sum_004+    tia_h_out_002_004+ sum_h_in_002_004- 260
Rh002_sum_004-    tia_h_out_002_004- sum_h_in_002_004+ 260
Rh002_sum_l_004   sum_h_in_002_004+ 0 650.0
Rh002_sum_fb_004  sum_h_in_002_004- sum_h_out_002_004 650.0
XUh002_sum_004    sum_h_in_002_004+ sum_h_in_002_004- Vcc+ Vcc- sum_h_out_002_004 MAX4223
* Neuron 5
Rh002_fb_005+     tia_h_in_002_005+ tia_h_out_002_005+ 4785.331062648607
Rh002_fb_005-     tia_h_in_002_005- tia_h_out_002_005- 4785.331062648607
XUh002_005+       0 tia_h_in_002_005+ Vcc+ Vcc- tia_h_out_002_005+ Ve OPA684_0
XUh002_005-       0 tia_h_in_002_005- Vcc+ Vcc- tia_h_out_002_005- Ve OPA684_0
Rh002_sum_005+    tia_h_out_002_005+ sum_h_in_002_005- 260
Rh002_sum_005-    tia_h_out_002_005- sum_h_in_002_005+ 260
Rh002_sum_l_005   sum_h_in_002_005+ 0 650.0
Rh002_sum_fb_005  sum_h_in_002_005- sum_h_out_002_005 650.0
XUh002_sum_005    sum_h_in_002_005+ sum_h_in_002_005- Vcc+ Vcc- sum_h_out_002_005 MAX4223
* Neuron 6
Rh002_fb_006+     tia_h_in_002_006+ tia_h_out_002_006+ 4785.331062648607
Rh002_fb_006-     tia_h_in_002_006- tia_h_out_002_006- 4785.331062648607
XUh002_006+       0 tia_h_in_002_006+ Vcc+ Vcc- tia_h_out_002_006+ Ve OPA684_0
XUh002_006-       0 tia_h_in_002_006- Vcc+ Vcc- tia_h_out_002_006- Ve OPA684_0
Rh002_sum_006+    tia_h_out_002_006+ sum_h_in_002_006- 260
Rh002_sum_006-    tia_h_out_002_006- sum_h_in_002_006+ 260
Rh002_sum_l_006   sum_h_in_002_006+ 0 650.0
Rh002_sum_fb_006  sum_h_in_002_006- sum_h_out_002_006 650.0
XUh002_sum_006    sum_h_in_002_006+ sum_h_in_002_006- Vcc+ Vcc- sum_h_out_002_006 MAX4223
* Neuron 7
Rh002_fb_007+     tia_h_in_002_007+ tia_h_out_002_007+ 4785.331062648607
Rh002_fb_007-     tia_h_in_002_007- tia_h_out_002_007- 4785.331062648607
XUh002_007+       0 tia_h_in_002_007+ Vcc+ Vcc- tia_h_out_002_007+ Ve OPA684_0
XUh002_007-       0 tia_h_in_002_007- Vcc+ Vcc- tia_h_out_002_007- Ve OPA684_0
Rh002_sum_007+    tia_h_out_002_007+ sum_h_in_002_007- 260
Rh002_sum_007-    tia_h_out_002_007- sum_h_in_002_007+ 260
Rh002_sum_l_007   sum_h_in_002_007+ 0 650.0
Rh002_sum_fb_007  sum_h_in_002_007- sum_h_out_002_007 650.0
XUh002_sum_007    sum_h_in_002_007+ sum_h_in_002_007- Vcc+ Vcc- sum_h_out_002_007 MAX4223
* Neuron 8
Rh002_fb_008+     tia_h_in_002_008+ tia_h_out_002_008+ 4785.331062648607
Rh002_fb_008-     tia_h_in_002_008- tia_h_out_002_008- 4785.331062648607
XUh002_008+       0 tia_h_in_002_008+ Vcc+ Vcc- tia_h_out_002_008+ Ve OPA684_0
XUh002_008-       0 tia_h_in_002_008- Vcc+ Vcc- tia_h_out_002_008- Ve OPA684_0
Rh002_sum_008+    tia_h_out_002_008+ sum_h_in_002_008- 260
Rh002_sum_008-    tia_h_out_002_008- sum_h_in_002_008+ 260
Rh002_sum_l_008   sum_h_in_002_008+ 0 650.0
Rh002_sum_fb_008  sum_h_in_002_008- sum_h_out_002_008 650.0
XUh002_sum_008    sum_h_in_002_008+ sum_h_in_002_008- Vcc+ Vcc- sum_h_out_002_008 MAX4223
* Neuron 9
Rh002_fb_009+     tia_h_in_002_009+ tia_h_out_002_009+ 4785.331062648607
Rh002_fb_009-     tia_h_in_002_009- tia_h_out_002_009- 4785.331062648607
XUh002_009+       0 tia_h_in_002_009+ Vcc+ Vcc- tia_h_out_002_009+ Ve OPA684_0
XUh002_009-       0 tia_h_in_002_009- Vcc+ Vcc- tia_h_out_002_009- Ve OPA684_0
Rh002_sum_009+    tia_h_out_002_009+ sum_h_in_002_009- 260
Rh002_sum_009-    tia_h_out_002_009- sum_h_in_002_009+ 260
Rh002_sum_l_009   sum_h_in_002_009+ 0 650.0
Rh002_sum_fb_009  sum_h_in_002_009- sum_h_out_002_009 650.0
XUh002_sum_009    sum_h_in_002_009+ sum_h_in_002_009- Vcc+ Vcc- sum_h_out_002_009 MAX4223
* Neuron 10
Rh002_fb_010+     tia_h_in_002_010+ tia_h_out_002_010+ 4785.331062648607
Rh002_fb_010-     tia_h_in_002_010- tia_h_out_002_010- 4785.331062648607
XUh002_010+       0 tia_h_in_002_010+ Vcc+ Vcc- tia_h_out_002_010+ Ve OPA684_0
XUh002_010-       0 tia_h_in_002_010- Vcc+ Vcc- tia_h_out_002_010- Ve OPA684_0
Rh002_sum_010+    tia_h_out_002_010+ sum_h_in_002_010- 260
Rh002_sum_010-    tia_h_out_002_010- sum_h_in_002_010+ 260
Rh002_sum_l_010   sum_h_in_002_010+ 0 650.0
Rh002_sum_fb_010  sum_h_in_002_010- sum_h_out_002_010 650.0
XUh002_sum_010    sum_h_in_002_010+ sum_h_in_002_010- Vcc+ Vcc- sum_h_out_002_010 MAX4223

* Layer 002
* Neuron 1
Rh003_fb_001+     tia_h_in_003_001+ tia_h_out_003_001+ 4785.331062648607
Rh003_fb_001-     tia_h_in_003_001- tia_h_out_003_001- 4785.331062648607
XUh003_001+       0 tia_h_in_003_001+ Vcc+ Vcc- tia_h_out_003_001+ Ve OPA684_0
XUh003_001-       0 tia_h_in_003_001- Vcc+ Vcc- tia_h_out_003_001- Ve OPA684_0
Rh003_sum_001+    tia_h_out_003_001+ sum_h_in_003_001- 260
Rh003_sum_001-    tia_h_out_003_001- sum_h_in_003_001+ 260
Rh003_sum_l_001   sum_h_in_003_001+ 0 650.0
Rh003_sum_fb_001  sum_h_in_003_001- sum_h_out_003_001 650.0
XUh003_sum_001    sum_h_in_003_001+ sum_h_in_003_001- Vcc+ Vcc- sum_h_out_003_001 MAX4223


* ----- Activation function Hard-Tanh)


* Layer 000
* Neuron 1
* XHardTanh_h001_001 sum_h_out_001_001 hidden_activ_out_h001_001 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_001 sum_h_out_001_001 hidden_activ_out_h001_001 ReLU
*XSigmoid_001_001 sum_h_out_001_001 hidden_activ_out_h001_001 RNN_Sigmoid3_HA
* Neuron 2
* XHardTanh_h001_002 sum_h_out_001_002 hidden_activ_out_h001_002 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_002 sum_h_out_001_002 hidden_activ_out_h001_002 ReLU
*XSigmoid_001_002 sum_h_out_001_002 hidden_activ_out_h001_002 RNN_Sigmoid3_HA
* Neuron 3
* XHardTanh_h001_003 sum_h_out_001_003 hidden_activ_out_h001_003 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_003 sum_h_out_001_003 hidden_activ_out_h001_003 ReLU
*XSigmoid_001_003 sum_h_out_001_003 hidden_activ_out_h001_003 RNN_Sigmoid3_HA
* Neuron 4
* XHardTanh_h001_004 sum_h_out_001_004 hidden_activ_out_h001_004 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_004 sum_h_out_001_004 hidden_activ_out_h001_004 ReLU
*XSigmoid_001_004 sum_h_out_001_004 hidden_activ_out_h001_004 RNN_Sigmoid3_HA
* Neuron 5
* XHardTanh_h001_005 sum_h_out_001_005 hidden_activ_out_h001_005 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_005 sum_h_out_001_005 hidden_activ_out_h001_005 ReLU
*XSigmoid_001_005 sum_h_out_001_005 hidden_activ_out_h001_005 RNN_Sigmoid3_HA
* Neuron 6
* XHardTanh_h001_006 sum_h_out_001_006 hidden_activ_out_h001_006 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_006 sum_h_out_001_006 hidden_activ_out_h001_006 ReLU
*XSigmoid_001_006 sum_h_out_001_006 hidden_activ_out_h001_006 RNN_Sigmoid3_HA
* Neuron 7
* XHardTanh_h001_007 sum_h_out_001_007 hidden_activ_out_h001_007 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_007 sum_h_out_001_007 hidden_activ_out_h001_007 ReLU
*XSigmoid_001_007 sum_h_out_001_007 hidden_activ_out_h001_007 RNN_Sigmoid3_HA
* Neuron 8
* XHardTanh_h001_008 sum_h_out_001_008 hidden_activ_out_h001_008 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_008 sum_h_out_001_008 hidden_activ_out_h001_008 ReLU
*XSigmoid_001_008 sum_h_out_001_008 hidden_activ_out_h001_008 RNN_Sigmoid3_HA
* Neuron 9
* XHardTanh_h001_009 sum_h_out_001_009 hidden_activ_out_h001_009 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_009 sum_h_out_001_009 hidden_activ_out_h001_009 ReLU
*XSigmoid_001_009 sum_h_out_001_009 hidden_activ_out_h001_009 RNN_Sigmoid3_HA
* Neuron 10
* XHardTanh_h001_010 sum_h_out_001_010 hidden_activ_out_h001_010 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_010 sum_h_out_001_010 hidden_activ_out_h001_010 ReLU
*XSigmoid_001_010 sum_h_out_001_010 hidden_activ_out_h001_010 RNN_Sigmoid3_HA
* Neuron 11
* XHardTanh_h001_011 sum_h_out_001_011 hidden_activ_out_h001_011 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_011 sum_h_out_001_011 hidden_activ_out_h001_011 ReLU
*XSigmoid_001_011 sum_h_out_001_011 hidden_activ_out_h001_011 RNN_Sigmoid3_HA
* Neuron 12
* XHardTanh_h001_012 sum_h_out_001_012 hidden_activ_out_h001_012 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_012 sum_h_out_001_012 hidden_activ_out_h001_012 ReLU
*XSigmoid_001_012 sum_h_out_001_012 hidden_activ_out_h001_012 RNN_Sigmoid3_HA
* Neuron 13
* XHardTanh_h001_013 sum_h_out_001_013 hidden_activ_out_h001_013 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_013 sum_h_out_001_013 hidden_activ_out_h001_013 ReLU
*XSigmoid_001_013 sum_h_out_001_013 hidden_activ_out_h001_013 RNN_Sigmoid3_HA
* Neuron 14
* XHardTanh_h001_014 sum_h_out_001_014 hidden_activ_out_h001_014 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_014 sum_h_out_001_014 hidden_activ_out_h001_014 ReLU
*XSigmoid_001_014 sum_h_out_001_014 hidden_activ_out_h001_014 RNN_Sigmoid3_HA
* Neuron 15
* XHardTanh_h001_015 sum_h_out_001_015 hidden_activ_out_h001_015 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_015 sum_h_out_001_015 hidden_activ_out_h001_015 ReLU
*XSigmoid_001_015 sum_h_out_001_015 hidden_activ_out_h001_015 RNN_Sigmoid3_HA
* Neuron 16
* XHardTanh_h001_016 sum_h_out_001_016 hidden_activ_out_h001_016 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_016 sum_h_out_001_016 hidden_activ_out_h001_016 ReLU
*XSigmoid_001_016 sum_h_out_001_016 hidden_activ_out_h001_016 RNN_Sigmoid3_HA
* Neuron 17
* XHardTanh_h001_017 sum_h_out_001_017 hidden_activ_out_h001_017 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_017 sum_h_out_001_017 hidden_activ_out_h001_017 ReLU
*XSigmoid_001_017 sum_h_out_001_017 hidden_activ_out_h001_017 RNN_Sigmoid3_HA
* Neuron 18
* XHardTanh_h001_018 sum_h_out_001_018 hidden_activ_out_h001_018 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_018 sum_h_out_001_018 hidden_activ_out_h001_018 ReLU
*XSigmoid_001_018 sum_h_out_001_018 hidden_activ_out_h001_018 RNN_Sigmoid3_HA
* Neuron 19
* XHardTanh_h001_019 sum_h_out_001_019 hidden_activ_out_h001_019 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_019 sum_h_out_001_019 hidden_activ_out_h001_019 ReLU
*XSigmoid_001_019 sum_h_out_001_019 hidden_activ_out_h001_019 RNN_Sigmoid3_HA
* Neuron 20
* XHardTanh_h001_020 sum_h_out_001_020 hidden_activ_out_h001_020 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_020 sum_h_out_001_020 hidden_activ_out_h001_020 ReLU
*XSigmoid_001_020 sum_h_out_001_020 hidden_activ_out_h001_020 RNN_Sigmoid3_HA

* Layer 001
* Neuron 1
* XHardTanh_h002_001 sum_h_out_002_001 hidden_activ_out_h002_001 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_001 sum_h_out_002_001 hidden_activ_out_h002_001 ReLU
*XSigmoid_002_001 sum_h_out_002_001 hidden_activ_out_h002_001 RNN_Sigmoid3_HA
* Neuron 2
* XHardTanh_h002_002 sum_h_out_002_002 hidden_activ_out_h002_002 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_002 sum_h_out_002_002 hidden_activ_out_h002_002 ReLU
*XSigmoid_002_002 sum_h_out_002_002 hidden_activ_out_h002_002 RNN_Sigmoid3_HA
* Neuron 3
* XHardTanh_h002_003 sum_h_out_002_003 hidden_activ_out_h002_003 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_003 sum_h_out_002_003 hidden_activ_out_h002_003 ReLU
*XSigmoid_002_003 sum_h_out_002_003 hidden_activ_out_h002_003 RNN_Sigmoid3_HA
* Neuron 4
* XHardTanh_h002_004 sum_h_out_002_004 hidden_activ_out_h002_004 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_004 sum_h_out_002_004 hidden_activ_out_h002_004 ReLU
*XSigmoid_002_004 sum_h_out_002_004 hidden_activ_out_h002_004 RNN_Sigmoid3_HA
* Neuron 5
* XHardTanh_h002_005 sum_h_out_002_005 hidden_activ_out_h002_005 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_005 sum_h_out_002_005 hidden_activ_out_h002_005 ReLU
*XSigmoid_002_005 sum_h_out_002_005 hidden_activ_out_h002_005 RNN_Sigmoid3_HA
* Neuron 6
* XHardTanh_h002_006 sum_h_out_002_006 hidden_activ_out_h002_006 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_006 sum_h_out_002_006 hidden_activ_out_h002_006 ReLU
*XSigmoid_002_006 sum_h_out_002_006 hidden_activ_out_h002_006 RNN_Sigmoid3_HA
* Neuron 7
* XHardTanh_h002_007 sum_h_out_002_007 hidden_activ_out_h002_007 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_007 sum_h_out_002_007 hidden_activ_out_h002_007 ReLU
*XSigmoid_002_007 sum_h_out_002_007 hidden_activ_out_h002_007 RNN_Sigmoid3_HA
* Neuron 8
* XHardTanh_h002_008 sum_h_out_002_008 hidden_activ_out_h002_008 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_008 sum_h_out_002_008 hidden_activ_out_h002_008 ReLU
*XSigmoid_002_008 sum_h_out_002_008 hidden_activ_out_h002_008 RNN_Sigmoid3_HA
* Neuron 9
* XHardTanh_h002_009 sum_h_out_002_009 hidden_activ_out_h002_009 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_009 sum_h_out_002_009 hidden_activ_out_h002_009 ReLU
*XSigmoid_002_009 sum_h_out_002_009 hidden_activ_out_h002_009 RNN_Sigmoid3_HA
* Neuron 10
* XHardTanh_h002_010 sum_h_out_002_010 hidden_activ_out_h002_010 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_010 sum_h_out_002_010 hidden_activ_out_h002_010 ReLU
*XSigmoid_002_010 sum_h_out_002_010 hidden_activ_out_h002_010 RNN_Sigmoid3_HA

* Layer 002
* Neuron 1
* XHardTanh_h003_001 sum_h_out_003_001 hidden_activ_out_h003_001 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_003_001 sum_h_out_003_001 hidden_activ_out_h003_001 ReLU
*XSigmoid_003_001 sum_h_out_003_001 hidden_activ_out_h003_001 RNN_Sigmoid3_HA


.END