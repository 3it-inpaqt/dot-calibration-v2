*
XX1 in out rnn_sigmoid3_ha
V1 in 0 PWL(0 -2 10u 2)

.print tran format=raw file=plot/Test_RNN_Sigmoid3_HA_xyce.raw v(*)
.tran 0 10u 10n
.include "..\models\180nm_bulk.txt"
.include "Sigmoid3_HA.spice"
.backanno
.end
nno
.end
