* Netlist that describe the physical circuit (components and connexions between them) to simulate, in Xyce formalism.
* To make the translation from any network size, the circuit is scaled up automatically using Jinja template engine.
*
* Xyce: https://xyce.sandia.gov
* Jinja: https://jinja.palletsprojects.com

* ======================== Simulation parameters ==========================

.TRAN 0.30ns 331.00ns

* OPTIONS TIMEINT change the time integration parameters
* ERROPTION (If 0 Local Truncation Error is used)
* METHOD: Time integration method
* NLMIN, NLMAX:  lower and upper bound for the desired number of nonlinear iterations
* DELMAX: The maximum time step-size used
* This additional line allows to fix convergence problem but increases the simulation time
* List variables to save in the result table
.PRINT TRAN V(sum_h_out_003_001) V(hidden_activ_out_h003_001)
+ V(i_001) V(i_002) V(i_003) V(i_004) V(i_005) V(i_006) V(i_007) V(i_008) V(i_009) V(i_010) V(i_011) V(i_012) V(i_013) V(i_014) V(i_015) V(i_016) V(i_017) V(i_018) V(i_019) V(i_020) V(i_021) V(i_022) V(i_023) V(i_024) V(i_025) V(i_026) V(i_027) V(i_028) V(i_029) V(i_030) V(i_031) V(i_032) V(i_033) V(i_034) V(i_035) V(i_036) V(i_037) V(i_038) V(i_039) V(i_040) V(i_041) V(i_042) V(i_043) V(i_044) V(i_045) V(i_046) V(i_047) V(i_048) V(i_049) V(i_050) V(i_051) V(i_052) V(i_053) V(i_054) V(i_055) V(i_056) V(i_057) V(i_058) V(i_059) V(i_060) V(i_061) V(i_062) V(i_063) V(i_064)
+ V(sum_h_out_001_001) V(hidden_activ_out_h001_001) V(sum_h_out_001_002) V(hidden_activ_out_h001_002) V(sum_h_out_001_003) V(hidden_activ_out_h001_003) V(sum_h_out_001_004) V(hidden_activ_out_h001_004) V(sum_h_out_001_005) V(hidden_activ_out_h001_005) V(sum_h_out_001_006) V(hidden_activ_out_h001_006) V(sum_h_out_001_007) V(hidden_activ_out_h001_007) V(sum_h_out_001_008) V(hidden_activ_out_h001_008) V(sum_h_out_001_009) V(hidden_activ_out_h001_009) V(sum_h_out_001_010) V(hidden_activ_out_h001_010) V(sum_h_out_001_011) V(hidden_activ_out_h001_011) V(sum_h_out_001_012) V(hidden_activ_out_h001_012) V(sum_h_out_001_013) V(hidden_activ_out_h001_013) V(sum_h_out_001_014) V(hidden_activ_out_h001_014) V(sum_h_out_001_015) V(hidden_activ_out_h001_015) V(sum_h_out_001_016) V(hidden_activ_out_h001_016) V(sum_h_out_001_017) V(hidden_activ_out_h001_017) V(sum_h_out_001_018) V(hidden_activ_out_h001_018) V(sum_h_out_001_019) V(hidden_activ_out_h001_019) V(sum_h_out_001_020) V(hidden_activ_out_h001_020)
+ V(tia_h_out_001_001+) V(tia_h_out_001_001-) V(tia_h_out_001_002+) V(tia_h_out_001_002-) V(tia_h_out_001_003+) V(tia_h_out_001_003-) V(tia_h_out_001_004+) V(tia_h_out_001_004-) V(tia_h_out_001_005+) V(tia_h_out_001_005-) V(tia_h_out_001_006+) V(tia_h_out_001_006-) V(tia_h_out_001_007+) V(tia_h_out_001_007-) V(tia_h_out_001_008+) V(tia_h_out_001_008-) V(tia_h_out_001_009+) V(tia_h_out_001_009-) V(tia_h_out_001_010+) V(tia_h_out_001_010-) V(tia_h_out_001_011+) V(tia_h_out_001_011-) V(tia_h_out_001_012+) V(tia_h_out_001_012-) V(tia_h_out_001_013+) V(tia_h_out_001_013-) V(tia_h_out_001_014+) V(tia_h_out_001_014-) V(tia_h_out_001_015+) V(tia_h_out_001_015-) V(tia_h_out_001_016+) V(tia_h_out_001_016-) V(tia_h_out_001_017+) V(tia_h_out_001_017-) V(tia_h_out_001_018+) V(tia_h_out_001_018-) V(tia_h_out_001_019+) V(tia_h_out_001_019-) V(tia_h_out_001_020+) V(tia_h_out_001_020-)
+ V(b_001)
+ V(sum_h_out_002_001) V(hidden_activ_out_h002_001) V(sum_h_out_002_002) V(hidden_activ_out_h002_002) V(sum_h_out_002_003) V(hidden_activ_out_h002_003) V(sum_h_out_002_004) V(hidden_activ_out_h002_004) V(sum_h_out_002_005) V(hidden_activ_out_h002_005) V(sum_h_out_002_006) V(hidden_activ_out_h002_006) V(sum_h_out_002_007) V(hidden_activ_out_h002_007) V(sum_h_out_002_008) V(hidden_activ_out_h002_008) V(sum_h_out_002_009) V(hidden_activ_out_h002_009) V(sum_h_out_002_010) V(hidden_activ_out_h002_010)
+ V(tia_h_out_002_001+) V(tia_h_out_002_001-) V(tia_h_out_002_002+) V(tia_h_out_002_002-) V(tia_h_out_002_003+) V(tia_h_out_002_003-) V(tia_h_out_002_004+) V(tia_h_out_002_004-) V(tia_h_out_002_005+) V(tia_h_out_002_005-) V(tia_h_out_002_006+) V(tia_h_out_002_006-) V(tia_h_out_002_007+) V(tia_h_out_002_007-) V(tia_h_out_002_008+) V(tia_h_out_002_008-) V(tia_h_out_002_009+) V(tia_h_out_002_009-) V(tia_h_out_002_010+) V(tia_h_out_002_010-)
+ V(b_002)
+ V(sum_h_out_003_001) V(hidden_activ_out_h003_001)
+ V(tia_h_out_003_001+) V(tia_h_out_003_001-)
+ V(b_003)

* =============================== Models ==================================

* Call the defined components model from the specified path
*.INCLUDE "./components/MAX4223.sub"
.INCLUDE "./components/TLV3501.sub"
*.INCLUDE "./components/OPA684.sub"

* Import custom sub-circuits
.INCLUDE "./components/activations.sub"
.INCLUDE "./components/lumped_line.sub"
.INCLUDE "./components/Sigmoid3_HA.spice"

* Define diode model
.MODEL D_BAV74_1 D( IS=2.073F N=1 BV=50 IBV=100N RS=1.336 
+      CJO=2P VJ=750M M=330M FC=500M TT=5.771N 
+      EG=1.11 XTI=3 KF=0 AF=1 )

* ============================== Voltages =================================

* ----- Input pulses
* Vi_num: The input voltage as pulse sequences
Vi_001    i_001    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.083V 300.00ns 1.083V 301.00ns 0.950V
Vi_002    i_002    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.035V 300.00ns 1.035V 301.00ns 0.950V
Vi_003    i_003    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.000V 300.00ns 1.000V 301.00ns 0.950V
Vi_004    i_004    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.972V 300.00ns 0.972V 301.00ns 0.950V
Vi_005    i_005    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.009V 300.00ns 1.009V 301.00ns 0.950V
Vi_006    i_006    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.995V 300.00ns 0.995V 301.00ns 0.950V
Vi_007    i_007    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.042V 300.00ns 1.042V 301.00ns 0.950V
Vi_008    i_008    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.950V 300.00ns 0.950V 301.00ns 0.950V
Vi_009    i_009    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.080V 300.00ns 1.080V 301.00ns 0.950V
Vi_010    i_010    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.039V 300.00ns 1.039V 301.00ns 0.950V
Vi_011    i_011    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.995V 300.00ns 0.995V 301.00ns 0.950V
Vi_012    i_012    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.005V 300.00ns 1.005V 301.00ns 0.950V
Vi_013    i_013    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.010V 300.00ns 1.010V 301.00ns 0.950V
Vi_014    i_014    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.038V 300.00ns 1.038V 301.00ns 0.950V
Vi_015    i_015    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.053V 300.00ns 1.053V 301.00ns 0.950V
Vi_016    i_016    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.960V 300.00ns 0.960V 301.00ns 0.950V
Vi_017    i_017    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.073V 300.00ns 1.073V 301.00ns 0.950V
Vi_018    i_018    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.050V 300.00ns 1.050V 301.00ns 0.950V
Vi_019    i_019    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.992V 300.00ns 0.992V 301.00ns 0.950V
Vi_020    i_020    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.025V 300.00ns 1.025V 301.00ns 0.950V
Vi_021    i_021    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.072V 300.00ns 1.072V 301.00ns 0.950V
Vi_022    i_022    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.035V 300.00ns 1.035V 301.00ns 0.950V
Vi_023    i_023    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.081V 300.00ns 1.081V 301.00ns 0.950V
Vi_024    i_024    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.996V 300.00ns 0.996V 301.00ns 0.950V
Vi_025    i_025    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.104V 300.00ns 1.104V 301.00ns 0.950V
Vi_026    i_026    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.054V 300.00ns 1.054V 301.00ns 0.950V
Vi_027    i_027    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.019V 300.00ns 1.019V 301.00ns 0.950V
Vi_028    i_028    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.028V 300.00ns 1.028V 301.00ns 0.950V
Vi_029    i_029    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.034V 300.00ns 1.034V 301.00ns 0.950V
Vi_030    i_030    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.049V 300.00ns 1.049V 301.00ns 0.950V
Vi_031    i_031    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.072V 300.00ns 1.072V 301.00ns 0.950V
Vi_032    i_032    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 0.995V 300.00ns 0.995V 301.00ns 0.950V
Vi_033    i_033    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.130V 300.00ns 1.130V 301.00ns 0.950V
Vi_034    i_034    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.073V 300.00ns 1.073V 301.00ns 0.950V
Vi_035    i_035    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.030V 300.00ns 1.030V 301.00ns 0.950V
Vi_036    i_036    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.023V 300.00ns 1.023V 301.00ns 0.950V
Vi_037    i_037    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.087V 300.00ns 1.087V 301.00ns 0.950V
Vi_038    i_038    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.066V 300.00ns 1.066V 301.00ns 0.950V
Vi_039    i_039    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.086V 300.00ns 1.086V 301.00ns 0.950V
Vi_040    i_040    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.019V 300.00ns 1.019V 301.00ns 0.950V
Vi_041    i_041    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.150V 300.00ns 1.150V 301.00ns 0.950V
Vi_042    i_042    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.091V 300.00ns 1.091V 301.00ns 0.950V
Vi_043    i_043    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.036V 300.00ns 1.036V 301.00ns 0.950V
Vi_044    i_044    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.042V 300.00ns 1.042V 301.00ns 0.950V
Vi_045    i_045    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.094V 300.00ns 1.094V 301.00ns 0.950V
Vi_046    i_046    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.075V 300.00ns 1.075V 301.00ns 0.950V
Vi_047    i_047    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.103V 300.00ns 1.103V 301.00ns 0.950V
Vi_048    i_048    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.023V 300.00ns 1.023V 301.00ns 0.950V
Vi_049    i_049    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.136V 300.00ns 1.136V 301.00ns 0.950V
Vi_050    i_050    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.109V 300.00ns 1.109V 301.00ns 0.950V
Vi_051    i_051    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.062V 300.00ns 1.062V 301.00ns 0.950V
Vi_052    i_052    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.044V 300.00ns 1.044V 301.00ns 0.950V
Vi_053    i_053    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.100V 300.00ns 1.100V 301.00ns 0.950V
Vi_054    i_054    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.085V 300.00ns 1.085V 301.00ns 0.950V
Vi_055    i_055    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.091V 300.00ns 1.091V 301.00ns 0.950V
Vi_056    i_056    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.020V 300.00ns 1.020V 301.00ns 0.950V
Vi_057    i_057    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.133V 300.00ns 1.133V 301.00ns 0.950V
Vi_058    i_058    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.107V 300.00ns 1.107V 301.00ns 0.950V
Vi_059    i_059    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.074V 300.00ns 1.074V 301.00ns 0.950V
Vi_060    i_060    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.045V 300.00ns 1.045V 301.00ns 0.950V
Vi_061    i_061    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.115V 300.00ns 1.115V 301.00ns 0.950V
Vi_062    i_062    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.057V 300.00ns 1.057V 301.00ns 0.950V
Vi_063    i_063    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.135V 300.00ns 1.135V 301.00ns 0.950V
Vi_064    i_064    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.033V 300.00ns 1.033V 301.00ns 0.950V

* Vb_num: The bias voltage as pulse sequences

Vb_001    b_001    0    PWL 0.00ns 0.950V 1.00ns 0.950V 2.00ns 1.150V 300.00ns 1.150V 301.00ns 0.950V
Vb_002    b_002    0    PWL 0.00ns 0.950V 11.00ns 0.950V 12.00ns 1.150V 310.00ns 1.150V 311.00ns 0.950V
Vb_003    b_003    0    PWL 0.00ns 0.950V 21.00ns 0.950V 22.00ns 1.150V 320.00ns 1.150V 321.00ns 0.950V

Ve        Ve       0    3
Vcc-      Vcc-     0    -5
Vcc+      Vcc+     0    5

* ============================ NN Parameters ==============================
* Parameters (weights and bias) naming convention: "Rl_i_j+" where:
*   R: Always "R" to inform Xyce it is a resistance
*   l: layer name, "h" for the hidden and output layers and "b" for the biases.
*   i: index of the weight of a neuron (start from 1)
*   j: index of the neuron (start from 1)
*   +: parameter polarity, + or -

* ----------------------------- Layers -----------------------------


* ----- Weights
* Layer 001

* Neuron 1
Rh001_001_001+    i_001    tia_h_in_001_001+    15128.645440125883
Rh001_001_001-    i_001    tia_h_in_001_001-    11474.80562712368
Rh001_002_001+    i_002    tia_h_in_001_001+    15087.564080154194
Rh001_002_001-    i_002    tia_h_in_001_001-    11026.319916672737
Rh001_003_001+    i_003    tia_h_in_001_001+    14847.548166584069
Rh001_003_001-    i_003    tia_h_in_001_001-    14870.883491042723
Rh001_004_001+    i_004    tia_h_in_001_001+    11565.267725398844
Rh001_004_001-    i_004    tia_h_in_001_001-    15108.430622479931
Rh001_005_001+    i_005    tia_h_in_001_001+    11021.394107780849
Rh001_005_001-    i_005    tia_h_in_001_001-    15022.787015131626
Rh001_006_001+    i_006    tia_h_in_001_001+    11711.942577320095
Rh001_006_001-    i_006    tia_h_in_001_001-    14991.586341827804
Rh001_007_001+    i_007    tia_h_in_001_001+    15150.05848069798
Rh001_007_001-    i_007    tia_h_in_001_001-    14276.855380459541
Rh001_008_001+    i_008    tia_h_in_001_001+    15116.854420638254
Rh001_008_001-    i_008    tia_h_in_001_001-    13612.848211238468
Rh001_009_001+    i_009    tia_h_in_001_001+    14989.464455914253
Rh001_009_001-    i_009    tia_h_in_001_001-    14250.32100331042
Rh001_010_001+    i_010    tia_h_in_001_001+    14101.172277728057
Rh001_010_001-    i_010    tia_h_in_001_001-    14975.12428797091
Rh001_011_001+    i_011    tia_h_in_001_001+    11965.079991118457
Rh001_011_001-    i_011    tia_h_in_001_001-    15069.739034413593
Rh001_012_001+    i_012    tia_h_in_001_001+    12806.157935707408
Rh001_012_001-    i_012    tia_h_in_001_001-    14797.290350669084
Rh001_013_001+    i_013    tia_h_in_001_001+    13485.666507664318
Rh001_013_001-    i_013    tia_h_in_001_001-    14876.993082012015
Rh001_014_001+    i_014    tia_h_in_001_001+    14949.688446712637
Rh001_014_001-    i_014    tia_h_in_001_001-    13618.269430368162
Rh001_015_001+    i_015    tia_h_in_001_001+    15013.486830013226
Rh001_015_001-    i_015    tia_h_in_001_001-    12110.276703066007
Rh001_016_001+    i_016    tia_h_in_001_001+    14911.73550663397
Rh001_016_001-    i_016    tia_h_in_001_001-    14262.36971425265
Rh001_017_001+    i_017    tia_h_in_001_001+    15151.34126685275
Rh001_017_001-    i_017    tia_h_in_001_001-    13681.128799180902
Rh001_018_001+    i_018    tia_h_in_001_001+    13006.029923655815
Rh001_018_001-    i_018    tia_h_in_001_001-    14877.62711116211
Rh001_019_001+    i_019    tia_h_in_001_001+    5000
Rh001_019_001-    i_019    tia_h_in_001_001-    5000
Rh001_020_001+    i_020    tia_h_in_001_001+    11650.936987687683
Rh001_020_001-    i_020    tia_h_in_001_001-    15219.636750997528
Rh001_021_001+    i_021    tia_h_in_001_001+    14375.617645413031
Rh001_021_001-    i_021    tia_h_in_001_001-    14759.77444020825
Rh001_022_001+    i_022    tia_h_in_001_001+    15074.72843672886
Rh001_022_001-    i_022    tia_h_in_001_001-    13752.761571248235
Rh001_023_001+    i_023    tia_h_in_001_001+    15040.2040179465
Rh001_023_001-    i_023    tia_h_in_001_001-    13833.312461969801
Rh001_024_001+    i_024    tia_h_in_001_001+    5000
Rh001_024_001-    i_024    tia_h_in_001_001-    12487.221183087697
Rh001_025_001+    i_025    tia_h_in_001_001+    12528.030587036585
Rh001_025_001-    i_025    tia_h_in_001_001-    15077.559334405898
Rh001_026_001+    i_026    tia_h_in_001_001+    13659.466093848629
Rh001_026_001-    i_026    tia_h_in_001_001-    15002.048156141673
Rh001_027_001+    i_027    tia_h_in_001_001+    11993.183931238904
Rh001_027_001-    i_027    tia_h_in_001_001-    5000
Rh001_028_001+    i_028    tia_h_in_001_001+    14630.71115150191
Rh001_028_001-    i_028    tia_h_in_001_001-    15147.81508315075
Rh001_029_001+    i_029    tia_h_in_001_001+    15145.90386474744
Rh001_029_001-    i_029    tia_h_in_001_001-    12849.891992043948
Rh001_030_001+    i_030    tia_h_in_001_001+    15094.430676044014
Rh001_030_001-    i_030    tia_h_in_001_001-    13275.766524532739
Rh001_031_001+    i_031    tia_h_in_001_001+    14873.931726607745
Rh001_031_001-    i_031    tia_h_in_001_001-    5000
Rh001_032_001+    i_032    tia_h_in_001_001+    14030.842697361802
Rh001_032_001-    i_032    tia_h_in_001_001-    15220.16565748861
Rh001_033_001+    i_033    tia_h_in_001_001+    5000
Rh001_033_001-    i_033    tia_h_in_001_001-    14900.15162491189
Rh001_034_001+    i_034    tia_h_in_001_001+    5000
Rh001_034_001-    i_034    tia_h_in_001_001-    14736.823832551387
Rh001_035_001+    i_035    tia_h_in_001_001+    14947.471000985364
Rh001_035_001-    i_035    tia_h_in_001_001-    14906.046983335713
Rh001_036_001+    i_036    tia_h_in_001_001+    14966.815413486076
Rh001_036_001-    i_036    tia_h_in_001_001-    14488.727163104022
Rh001_037_001+    i_037    tia_h_in_001_001+    14884.980723576462
Rh001_037_001-    i_037    tia_h_in_001_001-    14493.73909477778
Rh001_038_001+    i_038    tia_h_in_001_001+    15214.11540653877
Rh001_038_001-    i_038    tia_h_in_001_001-    5000
Rh001_039_001+    i_039    tia_h_in_001_001+    15090.60904728418
Rh001_039_001-    i_039    tia_h_in_001_001-    14050.615034001908
Rh001_040_001+    i_040    tia_h_in_001_001+    13665.01478020349
Rh001_040_001-    i_040    tia_h_in_001_001-    14735.446279437061
Rh001_041_001+    i_041    tia_h_in_001_001+    13376.103860585206
Rh001_041_001-    i_041    tia_h_in_001_001-    15050.570225968273
Rh001_042_001+    i_042    tia_h_in_001_001+    15102.394419059468
Rh001_042_001-    i_042    tia_h_in_001_001-    13941.573472860382
Rh001_043_001+    i_043    tia_h_in_001_001+    15135.614889441
Rh001_043_001-    i_043    tia_h_in_001_001-    15167.75069257208
Rh001_044_001+    i_044    tia_h_in_001_001+    15092.86975970757
Rh001_044_001-    i_044    tia_h_in_001_001-    15000
Rh001_045_001+    i_045    tia_h_in_001_001+    14964.447073298023
Rh001_045_001-    i_045    tia_h_in_001_001-    13745.319250098542
Rh001_046_001+    i_046    tia_h_in_001_001+    14925.203582027936
Rh001_046_001-    i_046    tia_h_in_001_001-    13621.258370255902
Rh001_047_001+    i_047    tia_h_in_001_001+    13808.977512270269
Rh001_047_001-    i_047    tia_h_in_001_001-    14923.455763230733
Rh001_048_001+    i_048    tia_h_in_001_001+    15000
Rh001_048_001-    i_048    tia_h_in_001_001-    15206.61630813718
Rh001_049_001+    i_049    tia_h_in_001_001+    13195.964356039802
Rh001_049_001-    i_049    tia_h_in_001_001-    15116.417439679839
Rh001_050_001+    i_050    tia_h_in_001_001+    13261.992238140856
Rh001_050_001-    i_050    tia_h_in_001_001-    15088.693154064662
Rh001_051_001+    i_051    tia_h_in_001_001+    15082.47152212622
Rh001_051_001-    i_051    tia_h_in_001_001-    14480.517528450198
Rh001_052_001+    i_052    tia_h_in_001_001+    15072.217048442244
Rh001_052_001-    i_052    tia_h_in_001_001-    13895.90763425265
Rh001_053_001+    i_053    tia_h_in_001_001+    14998.350244808273
Rh001_053_001-    i_053    tia_h_in_001_001-    13043.618512432366
Rh001_054_001+    i_054    tia_h_in_001_001+    15143.41283007239
Rh001_054_001-    i_054    tia_h_in_001_001-    5000
Rh001_055_001+    i_055    tia_h_in_001_001+    14215.580765570108
Rh001_055_001-    i_055    tia_h_in_001_001-    14995.397031051358
Rh001_056_001+    i_056    tia_h_in_001_001+    14903.719507046917
Rh001_056_001-    i_056    tia_h_in_001_001-    13653.47609174428
Rh001_057_001+    i_057    tia_h_in_001_001+    5000
Rh001_057_001-    i_057    tia_h_in_001_001-    15109.244136594276
Rh001_058_001+    i_058    tia_h_in_001_001+    15072.888588347781
Rh001_058_001-    i_058    tia_h_in_001_001-    14237.09442482208
Rh001_059_001+    i_059    tia_h_in_001_001+    15148.264708190763
Rh001_059_001-    i_059    tia_h_in_001_001-    10746.063733299425
Rh001_060_001+    i_060    tia_h_in_001_001+    15000
Rh001_060_001-    i_060    tia_h_in_001_001-    10881.016471736744
Rh001_061_001+    i_061    tia_h_in_001_001+    15066.093848303766
Rh001_061_001-    i_061    tia_h_in_001_001-    14772.525186942614
Rh001_062_001+    i_062    tia_h_in_001_001+    12862.380909640671
Rh001_062_001-    i_062    tia_h_in_001_001-    15282.22216474602
Rh001_063_001+    i_063    tia_h_in_001_001+    11679.44856263123
Rh001_063_001-    i_063    tia_h_in_001_001-    15058.73945461571
Rh001_064_001+    i_064    tia_h_in_001_001+    12289.079392465977
Rh001_064_001-    i_064    tia_h_in_001_001-    14987.198785999297

* Neuron 2
Rh001_001_002+    i_001    tia_h_in_001_002+    15014.858192219417
Rh001_001_002-    i_001    tia_h_in_001_002-    12126.496304319602
Rh001_002_002+    i_002    tia_h_in_001_002+    14991.318063416127
Rh001_002_002-    i_002    tia_h_in_001_002-    11637.842455905067
Rh001_003_002+    i_003    tia_h_in_001_002+    14987.747211368232
Rh001_003_002-    i_003    tia_h_in_001_002-    13666.477054581774
Rh001_004_002+    i_004    tia_h_in_001_002+    15162.76266218755
Rh001_004_002-    i_004    tia_h_in_001_002-    5000
Rh001_005_002+    i_005    tia_h_in_001_002+    14699.51086309548
Rh001_005_002-    i_005    tia_h_in_001_002-    13882.080271948676
Rh001_006_002+    i_006    tia_h_in_001_002+    14863.53849280884
Rh001_006_002-    i_006    tia_h_in_001_002-    12176.636677049293
Rh001_007_002+    i_007    tia_h_in_001_002+    15022.772945827308
Rh001_007_002-    i_007    tia_h_in_001_002-    11911.92633101433
Rh001_008_002+    i_008    tia_h_in_001_002+    15018.376557614129
Rh001_008_002-    i_008    tia_h_in_001_002-    12313.320438918636
Rh001_009_002+    i_009    tia_h_in_001_002+    15167.934208435043
Rh001_009_002-    i_009    tia_h_in_001_002-    11566.516393733944
Rh001_010_002+    i_010    tia_h_in_001_002+    13082.446815243347
Rh001_010_002-    i_010    tia_h_in_001_002-    15000
Rh001_011_002+    i_011    tia_h_in_001_002+    14978.330214835734
Rh001_011_002-    i_011    tia_h_in_001_002-    14355.696420576714
Rh001_012_002+    i_012    tia_h_in_001_002+    12849.671959331685
Rh001_012_002-    i_012    tia_h_in_001_002-    15208.860834281606
Rh001_013_002+    i_013    tia_h_in_001_002+    14996.02224595237
Rh001_013_002-    i_013    tia_h_in_001_002-    15058.441194482279
Rh001_014_002+    i_014    tia_h_in_001_002+    14905.389168083058
Rh001_014_002-    i_014    tia_h_in_001_002-    14796.512424366641
Rh001_015_002+    i_015    tia_h_in_001_002+    13635.629019265978
Rh001_015_002-    i_015    tia_h_in_001_002-    14876.229420071202
Rh001_016_002+    i_016    tia_h_in_001_002+    13821.258579435
Rh001_016_002-    i_016    tia_h_in_001_002-    15073.769492264326
Rh001_017_002+    i_017    tia_h_in_001_002+    12066.785123181895
Rh001_017_002-    i_017    tia_h_in_001_002-    15128.023865515574
Rh001_018_002+    i_018    tia_h_in_001_002+    14854.499887605054
Rh001_018_002-    i_018    tia_h_in_001_002-    5000
Rh001_019_002+    i_019    tia_h_in_001_002+    14901.048769737845
Rh001_019_002-    i_019    tia_h_in_001_002-    14987.227127706949
Rh001_020_002+    i_020    tia_h_in_001_002+    14948.10978570103
Rh001_020_002-    i_020    tia_h_in_001_002-    13919.268599267372
Rh001_021_002+    i_021    tia_h_in_001_002+    14506.784660528214
Rh001_021_002-    i_021    tia_h_in_001_002-    5000
Rh001_022_002+    i_022    tia_h_in_001_002+    12613.27985430457
Rh001_022_002-    i_022    tia_h_in_001_002-    14988.054536663536
Rh001_023_002+    i_023    tia_h_in_001_002+    11554.39524681432
Rh001_023_002-    i_023    tia_h_in_001_002-    14984.585239206472
Rh001_024_002+    i_024    tia_h_in_001_002+    11412.733545391617
Rh001_024_002-    i_024    tia_h_in_001_002-    15053.927930782094
Rh001_025_002+    i_025    tia_h_in_001_002+    13526.939491278996
Rh001_025_002-    i_025    tia_h_in_001_002-    5000
Rh001_026_002+    i_026    tia_h_in_001_002+    13442.669578375362
Rh001_026_002-    i_026    tia_h_in_001_002-    15188.31823845389
Rh001_027_002+    i_027    tia_h_in_001_002+    15095.289630394307
Rh001_027_002-    i_027    tia_h_in_001_002-    13775.12823909812
Rh001_028_002+    i_028    tia_h_in_001_002+    15120.017062423967
Rh001_028_002-    i_028    tia_h_in_001_002-    13390.361561875783
Rh001_029_002+    i_029    tia_h_in_001_002+    12668.614670918416
Rh001_029_002-    i_029    tia_h_in_001_002-    15116.339511185673
Rh001_030_002+    i_030    tia_h_in_001_002+    14340.76338793553
Rh001_030_002-    i_030    tia_h_in_001_002-    15239.989823537922
Rh001_031_002+    i_031    tia_h_in_001_002+    14502.349637492818
Rh001_031_002-    i_031    tia_h_in_001_002-    15171.567216095571
Rh001_032_002+    i_032    tia_h_in_001_002+    14920.43511304739
Rh001_032_002-    i_032    tia_h_in_001_002-    14872.324959608455
Rh001_033_002+    i_033    tia_h_in_001_002+    5000
Rh001_033_002-    i_033    tia_h_in_001_002-    14917.195326818915
Rh001_034_002+    i_034    tia_h_in_001_002+    13557.363196457249
Rh001_034_002-    i_034    tia_h_in_001_002-    5000
Rh001_035_002+    i_035    tia_h_in_001_002+    14682.918559356682
Rh001_035_002-    i_035    tia_h_in_001_002-    15035.509524014768
Rh001_036_002+    i_036    tia_h_in_001_002+    14972.408000606494
Rh001_036_002-    i_036    tia_h_in_001_002-    14295.712556326109
Rh001_037_002+    i_037    tia_h_in_001_002+    14586.115708109603
Rh001_037_002-    i_037    tia_h_in_001_002-    14938.492314747002
Rh001_038_002+    i_038    tia_h_in_001_002+    15020.476314478
Rh001_038_002-    i_038    tia_h_in_001_002-    14213.885040225727
Rh001_039_002+    i_039    tia_h_in_001_002+    15000
Rh001_039_002-    i_039    tia_h_in_001_002-    12520.315916128033
Rh001_040_002+    i_040    tia_h_in_001_002+    14920.108117004804
Rh001_040_002-    i_040    tia_h_in_001_002-    13548.188535574118
Rh001_041_002+    i_041    tia_h_in_001_002+    14804.362718359087
Rh001_041_002-    i_041    tia_h_in_001_002-    14944.118401083291
Rh001_042_002+    i_042    tia_h_in_001_002+    13831.653740869191
Rh001_042_002-    i_042    tia_h_in_001_002-    14930.95045613838
Rh001_043_002+    i_043    tia_h_in_001_002+    12187.741446146565
Rh001_043_002-    i_043    tia_h_in_001_002-    14836.667046562847
Rh001_044_002+    i_044    tia_h_in_001_002+    13602.082433355688
Rh001_044_002-    i_044    tia_h_in_001_002-    14994.550440262303
Rh001_045_002+    i_045    tia_h_in_001_002+    15354.523782738668
Rh001_045_002-    i_045    tia_h_in_001_002-    12773.016986278612
Rh001_046_002+    i_046    tia_h_in_001_002+    15087.690831523341
Rh001_046_002-    i_046    tia_h_in_001_002-    12626.885505128741
Rh001_047_002+    i_047    tia_h_in_001_002+    15094.401725930327
Rh001_047_002-    i_047    tia_h_in_001_002-    14420.534653498571
Rh001_048_002+    i_048    tia_h_in_001_002+    15084.169336209367
Rh001_048_002-    i_048    tia_h_in_001_002-    14370.571729512176
Rh001_049_002+    i_049    tia_h_in_001_002+    14833.706873248217
Rh001_049_002-    i_049    tia_h_in_001_002-    13359.690823896284
Rh001_050_002+    i_050    tia_h_in_001_002+    14740.784257417803
Rh001_050_002-    i_050    tia_h_in_001_002-    14715.34949338883
Rh001_051_002+    i_051    tia_h_in_001_002+    14847.05496460694
Rh001_051_002-    i_051    tia_h_in_001_002-    14591.900316128804
Rh001_052_002+    i_052    tia_h_in_001_002+    15008.018140592527
Rh001_052_002-    i_052    tia_h_in_001_002-    14548.440247521181
Rh001_053_002+    i_053    tia_h_in_001_002+    15190.407256812534
Rh001_053_002-    i_053    tia_h_in_001_002-    14284.901389356251
Rh001_054_002+    i_054    tia_h_in_001_002+    13510.9458473471
Rh001_054_002-    i_054    tia_h_in_001_002-    14908.84979399672
Rh001_055_002+    i_055    tia_h_in_001_002+    15000
Rh001_055_002-    i_055    tia_h_in_001_002-    13852.09260841928
Rh001_056_002+    i_056    tia_h_in_001_002+    15072.169328023983
Rh001_056_002-    i_056    tia_h_in_001_002-    15000
Rh001_057_002+    i_057    tia_h_in_001_002+    15256.575947650308
Rh001_057_002-    i_057    tia_h_in_001_002-    5000
Rh001_058_002+    i_058    tia_h_in_001_002+    15137.369367025945
Rh001_058_002-    i_058    tia_h_in_001_002-    14706.041578519995
Rh001_059_002+    i_059    tia_h_in_001_002+    15032.21913200211
Rh001_059_002-    i_059    tia_h_in_001_002-    13657.584688679288
Rh001_060_002+    i_060    tia_h_in_001_002+    15121.126069516595
Rh001_060_002-    i_060    tia_h_in_001_002-    14817.644424702661
Rh001_061_002+    i_061    tia_h_in_001_002+    15000
Rh001_061_002-    i_061    tia_h_in_001_002-    14979.674745518361
Rh001_062_002+    i_062    tia_h_in_001_002+    14201.303050220697
Rh001_062_002-    i_062    tia_h_in_001_002-    14927.950779007011
Rh001_063_002+    i_063    tia_h_in_001_002+    5000
Rh001_063_002-    i_063    tia_h_in_001_002-    14930.815935304096
Rh001_064_002+    i_064    tia_h_in_001_002+    14884.198715087072
Rh001_064_002-    i_064    tia_h_in_001_002-    13574.274494077936

* Neuron 3
Rh001_001_003+    i_001    tia_h_in_001_003+    15160.223754163213
Rh001_001_003-    i_001    tia_h_in_001_003-    13453.20300137503
Rh001_002_003+    i_002    tia_h_in_001_003+    15105.632922417093
Rh001_002_003-    i_002    tia_h_in_001_003-    13744.157244365853
Rh001_003_003+    i_003    tia_h_in_001_003+    11700.34439472623
Rh001_003_003-    i_003    tia_h_in_001_003-    14987.239306414864
Rh001_004_003+    i_004    tia_h_in_001_003+    10134.40251030774
Rh001_004_003-    i_004    tia_h_in_001_003-    15100.633534511953
Rh001_005_003+    i_005    tia_h_in_001_003+    12336.787312170753
Rh001_005_003-    i_005    tia_h_in_001_003-    15018.568934160614
Rh001_006_003+    i_006    tia_h_in_001_003+    14776.367557735704
Rh001_006_003-    i_006    tia_h_in_001_003-    14263.305197821228
Rh001_007_003+    i_007    tia_h_in_001_003+    15041.484395297854
Rh001_007_003-    i_007    tia_h_in_001_003-    12986.475297122615
Rh001_008_003+    i_008    tia_h_in_001_003+    15000
Rh001_008_003-    i_008    tia_h_in_001_003-    10703.589014343255
Rh001_009_003+    i_009    tia_h_in_001_003+    15000
Rh001_009_003-    i_009    tia_h_in_001_003-    14905.052593555329
Rh001_010_003+    i_010    tia_h_in_001_003+    13353.544404705643
Rh001_010_003-    i_010    tia_h_in_001_003-    15146.637525742342
Rh001_011_003+    i_011    tia_h_in_001_003+    12902.762679119009
Rh001_011_003-    i_011    tia_h_in_001_003-    15011.006426444708
Rh001_012_003+    i_012    tia_h_in_001_003+    15142.433838203644
Rh001_012_003-    i_012    tia_h_in_001_003-    14154.529424034059
Rh001_013_003+    i_013    tia_h_in_001_003+    5000
Rh001_013_003-    i_013    tia_h_in_001_003-    14889.72081441767
Rh001_014_003+    i_014    tia_h_in_001_003+    14824.096463892321
Rh001_014_003-    i_014    tia_h_in_001_003-    13422.332985767187
Rh001_015_003+    i_015    tia_h_in_001_003+    14806.892017852218
Rh001_015_003-    i_015    tia_h_in_001_003-    13190.492920238923
Rh001_016_003+    i_016    tia_h_in_001_003+    14946.001843668293
Rh001_016_003-    i_016    tia_h_in_001_003-    14306.51183666826
Rh001_017_003+    i_017    tia_h_in_001_003+    14303.301411410228
Rh001_017_003-    i_017    tia_h_in_001_003-    15069.216990691542
Rh001_018_003+    i_018    tia_h_in_001_003+    13784.52035568493
Rh001_018_003-    i_018    tia_h_in_001_003-    14998.234946509356
Rh001_019_003+    i_019    tia_h_in_001_003+    12098.663079530532
Rh001_019_003-    i_019    tia_h_in_001_003-    15106.893559476219
Rh001_020_003+    i_020    tia_h_in_001_003+    14335.565550363655
Rh001_020_003-    i_020    tia_h_in_001_003-    15154.524275279424
Rh001_021_003+    i_021    tia_h_in_001_003+    15031.920969308016
Rh001_021_003-    i_021    tia_h_in_001_003-    15004.979233757833
Rh001_022_003+    i_022    tia_h_in_001_003+    15056.041141189358
Rh001_022_003-    i_022    tia_h_in_001_003-    13197.56048955136
Rh001_023_003+    i_023    tia_h_in_001_003+    15246.02313846685
Rh001_023_003-    i_023    tia_h_in_001_003-    13519.34283152145
Rh001_024_003+    i_024    tia_h_in_001_003+    14779.88317935996
Rh001_024_003-    i_024    tia_h_in_001_003-    13668.207579308548
Rh001_025_003+    i_025    tia_h_in_001_003+    12603.372135348585
Rh001_025_003-    i_025    tia_h_in_001_003-    14966.7933602713
Rh001_026_003+    i_026    tia_h_in_001_003+    13659.694888980597
Rh001_026_003-    i_026    tia_h_in_001_003-    15024.633649906913
Rh001_027_003+    i_027    tia_h_in_001_003+    14216.616983505155
Rh001_027_003-    i_027    tia_h_in_001_003-    15188.082914982535
Rh001_028_003+    i_028    tia_h_in_001_003+    14971.991100758169
Rh001_028_003-    i_028    tia_h_in_001_003-    12980.887597104447
Rh001_029_003+    i_029    tia_h_in_001_003+    15004.403958644376
Rh001_029_003-    i_029    tia_h_in_001_003-    14262.589571678243
Rh001_030_003+    i_030    tia_h_in_001_003+    14952.590282756177
Rh001_030_003-    i_030    tia_h_in_001_003-    14258.687222370823
Rh001_031_003+    i_031    tia_h_in_001_003+    14448.431890894663
Rh001_031_003-    i_031    tia_h_in_001_003-    15115.154575756625
Rh001_032_003+    i_032    tia_h_in_001_003+    14102.438611567577
Rh001_032_003-    i_032    tia_h_in_001_003-    14838.276055935767
Rh001_033_003+    i_033    tia_h_in_001_003+    13460.736740889713
Rh001_033_003-    i_033    tia_h_in_001_003-    14987.202529068589
Rh001_034_003+    i_034    tia_h_in_001_003+    15000
Rh001_034_003-    i_034    tia_h_in_001_003-    14805.747953419876
Rh001_035_003+    i_035    tia_h_in_001_003+    14986.571759588527
Rh001_035_003-    i_035    tia_h_in_001_003-    12900.419220801787
Rh001_036_003+    i_036    tia_h_in_001_003+    5000
Rh001_036_003-    i_036    tia_h_in_001_003-    13808.196132667319
Rh001_037_003+    i_037    tia_h_in_001_003+    15101.265309169477
Rh001_037_003-    i_037    tia_h_in_001_003-    14412.910894065806
Rh001_038_003+    i_038    tia_h_in_001_003+    15087.415939508512
Rh001_038_003-    i_038    tia_h_in_001_003-    13639.572605387899
Rh001_039_003+    i_039    tia_h_in_001_003+    14696.443394926164
Rh001_039_003-    i_039    tia_h_in_001_003-    15128.460075640334
Rh001_040_003+    i_040    tia_h_in_001_003+    12172.485988680037
Rh001_040_003-    i_040    tia_h_in_001_003-    15053.90603909982
Rh001_041_003+    i_041    tia_h_in_001_003+    14531.370060730482
Rh001_041_003-    i_041    tia_h_in_001_003-    15113.722362300634
Rh001_042_003+    i_042    tia_h_in_001_003+    14922.591630544403
Rh001_042_003-    i_042    tia_h_in_001_003-    14875.129626645261
Rh001_043_003+    i_043    tia_h_in_001_003+    14923.744524323192
Rh001_043_003-    i_043    tia_h_in_001_003-    13113.273814698912
Rh001_044_003+    i_044    tia_h_in_001_003+    14950.717827953193
Rh001_044_003-    i_044    tia_h_in_001_003-    14402.976780045023
Rh001_045_003+    i_045    tia_h_in_001_003+    14936.812353922174
Rh001_045_003-    i_045    tia_h_in_001_003-    14454.120827228102
Rh001_046_003+    i_046    tia_h_in_001_003+    14459.093257939357
Rh001_046_003-    i_046    tia_h_in_001_003-    15074.318658056392
Rh001_047_003+    i_047    tia_h_in_001_003+    12032.233530969026
Rh001_047_003-    i_047    tia_h_in_001_003-    15088.095942313952
Rh001_048_003+    i_048    tia_h_in_001_003+    12189.978852385564
Rh001_048_003-    i_048    tia_h_in_001_003-    15103.00902734843
Rh001_049_003+    i_049    tia_h_in_001_003+    14386.347171621386
Rh001_049_003-    i_049    tia_h_in_001_003-    15029.056251359982
Rh001_050_003+    i_050    tia_h_in_001_003+    14777.42941957989
Rh001_050_003-    i_050    tia_h_in_001_003-    15000
Rh001_051_003+    i_051    tia_h_in_001_003+    14807.251315639232
Rh001_051_003-    i_051    tia_h_in_001_003-    14567.723650300619
Rh001_052_003+    i_052    tia_h_in_001_003+    14864.773580563822
Rh001_052_003-    i_052    tia_h_in_001_003-    13806.13925553174
Rh001_053_003+    i_053    tia_h_in_001_003+    15011.24146318223
Rh001_053_003-    i_053    tia_h_in_001_003-    13142.07674078023
Rh001_054_003+    i_054    tia_h_in_001_003+    15181.25042818565
Rh001_054_003-    i_054    tia_h_in_001_003-    14242.658208843608
Rh001_055_003+    i_055    tia_h_in_001_003+    12779.739366040327
Rh001_055_003-    i_055    tia_h_in_001_003-    15186.60453722753
Rh001_056_003+    i_056    tia_h_in_001_003+    14027.88060638031
Rh001_056_003-    i_056    tia_h_in_001_003-    15032.009046942601
Rh001_057_003+    i_057    tia_h_in_001_003+    15108.553929204685
Rh001_057_003-    i_057    tia_h_in_001_003-    12376.731393824879
Rh001_058_003+    i_058    tia_h_in_001_003+    15078.407280252502
Rh001_058_003-    i_058    tia_h_in_001_003-    13130.435491466777
Rh001_059_003+    i_059    tia_h_in_001_003+    15000
Rh001_059_003-    i_059    tia_h_in_001_003-    12097.874522421065
Rh001_060_003+    i_060    tia_h_in_001_003+    15196.299052344442
Rh001_060_003-    i_060    tia_h_in_001_003-    15000
Rh001_061_003+    i_061    tia_h_in_001_003+    13442.717453757206
Rh001_061_003-    i_061    tia_h_in_001_003-    5000
Rh001_062_003+    i_062    tia_h_in_001_003+    10487.540158442976
Rh001_062_003-    i_062    tia_h_in_001_003-    15075.226039094692
Rh001_063_003+    i_063    tia_h_in_001_003+    13341.579370068162
Rh001_063_003-    i_063    tia_h_in_001_003-    14921.32146491431
Rh001_064_003+    i_064    tia_h_in_001_003+    14197.886624969246
Rh001_064_003-    i_064    tia_h_in_001_003-    15053.386235375354

* Neuron 4
Rh001_001_004+    i_001    tia_h_in_001_004+    14823.085863592592
Rh001_001_004-    i_001    tia_h_in_001_004-    5000
Rh001_002_004+    i_002    tia_h_in_001_004+    15067.629293187143
Rh001_002_004-    i_002    tia_h_in_001_004-    14794.166036002895
Rh001_003_004+    i_003    tia_h_in_001_004+    5000
Rh001_003_004-    i_003    tia_h_in_001_004-    14900.264557483382
Rh001_004_004+    i_004    tia_h_in_001_004+    14598.228744824366
Rh001_004_004-    i_004    tia_h_in_001_004-    14957.593910094856
Rh001_005_004+    i_005    tia_h_in_001_004+    14931.778667230416
Rh001_005_004-    i_005    tia_h_in_001_004-    13508.238562385759
Rh001_006_004+    i_006    tia_h_in_001_004+    14862.618383681953
Rh001_006_004-    i_006    tia_h_in_001_004-    14486.788513683743
Rh001_007_004+    i_007    tia_h_in_001_004+    13689.65290039666
Rh001_007_004-    i_007    tia_h_in_001_004-    15142.331230228492
Rh001_008_004+    i_008    tia_h_in_001_004+    14475.663260322724
Rh001_008_004-    i_008    tia_h_in_001_004-    14806.700063622191
Rh001_009_004+    i_009    tia_h_in_001_004+    14947.225966144917
Rh001_009_004-    i_009    tia_h_in_001_004-    14912.004362744909
Rh001_010_004+    i_010    tia_h_in_001_004+    14836.47529127979
Rh001_010_004-    i_010    tia_h_in_001_004-    13938.468848195453
Rh001_011_004+    i_011    tia_h_in_001_004+    15096.923700169124
Rh001_011_004-    i_011    tia_h_in_001_004-    14045.3272787273
Rh001_012_004+    i_012    tia_h_in_001_004+    14995.246770950658
Rh001_012_004-    i_012    tia_h_in_001_004-    13716.611857906253
Rh001_013_004+    i_013    tia_h_in_001_004+    14970.219663940316
Rh001_013_004-    i_013    tia_h_in_001_004-    14427.85431734345
Rh001_014_004+    i_014    tia_h_in_001_004+    14613.062490291468
Rh001_014_004-    i_014    tia_h_in_001_004-    14826.518745024845
Rh001_015_004+    i_015    tia_h_in_001_004+    14146.71236792767
Rh001_015_004-    i_015    tia_h_in_001_004-    14889.351970717902
Rh001_016_004+    i_016    tia_h_in_001_004+    14421.633640143838
Rh001_016_004-    i_016    tia_h_in_001_004-    14827.901706152565
Rh001_017_004+    i_017    tia_h_in_001_004+    15211.640703231025
Rh001_017_004-    i_017    tia_h_in_001_004-    13598.067305624274
Rh001_018_004+    i_018    tia_h_in_001_004+    15039.773489967776
Rh001_018_004-    i_018    tia_h_in_001_004-    13936.318687523242
Rh001_019_004+    i_019    tia_h_in_001_004+    14894.635179901754
Rh001_019_004-    i_019    tia_h_in_001_004-    5000
Rh001_020_004+    i_020    tia_h_in_001_004+    13576.221798592536
Rh001_020_004-    i_020    tia_h_in_001_004-    15000
Rh001_021_004+    i_021    tia_h_in_001_004+    14754.511254803516
Rh001_021_004-    i_021    tia_h_in_001_004-    14979.342350295654
Rh001_022_004+    i_022    tia_h_in_001_004+    14984.05279343635
Rh001_022_004-    i_022    tia_h_in_001_004-    14257.796368079104
Rh001_023_004+    i_023    tia_h_in_001_004+    14442.336861961117
Rh001_023_004-    i_023    tia_h_in_001_004-    14996.616091331005
Rh001_024_004+    i_024    tia_h_in_001_004+    14973.985097585048
Rh001_024_004-    i_024    tia_h_in_001_004-    14132.903857212761
Rh001_025_004+    i_025    tia_h_in_001_004+    14921.333420355206
Rh001_025_004-    i_025    tia_h_in_001_004-    13883.215803381516
Rh001_026_004+    i_026    tia_h_in_001_004+    13874.226748535642
Rh001_026_004-    i_026    tia_h_in_001_004-    14935.577456994422
Rh001_027_004+    i_027    tia_h_in_001_004+    14900.98228554168
Rh001_027_004-    i_027    tia_h_in_001_004-    14276.493596737548
Rh001_028_004+    i_028    tia_h_in_001_004+    15147.310955854902
Rh001_028_004-    i_028    tia_h_in_001_004-    14607.303360562924
Rh001_029_004+    i_029    tia_h_in_001_004+    14882.846964453647
Rh001_029_004-    i_029    tia_h_in_001_004-    13472.509245778807
Rh001_030_004+    i_030    tia_h_in_001_004+    5000
Rh001_030_004-    i_030    tia_h_in_001_004-    14960.626285374961
Rh001_031_004+    i_031    tia_h_in_001_004+    13967.559227704533
Rh001_031_004-    i_031    tia_h_in_001_004-    15194.98003951113
Rh001_032_004+    i_032    tia_h_in_001_004+    14388.748747981486
Rh001_032_004-    i_032    tia_h_in_001_004-    14951.725938159729
Rh001_033_004+    i_033    tia_h_in_001_004+    15028.044325074092
Rh001_033_004-    i_033    tia_h_in_001_004-    13807.212894195989
Rh001_034_004+    i_034    tia_h_in_001_004+    15020.266927234623
Rh001_034_004-    i_034    tia_h_in_001_004-    13447.403764380417
Rh001_035_004+    i_035    tia_h_in_001_004+    14907.323832126545
Rh001_035_004-    i_035    tia_h_in_001_004-    13906.957875727516
Rh001_036_004+    i_036    tia_h_in_001_004+    14148.99288709543
Rh001_036_004-    i_036    tia_h_in_001_004-    15212.476358893267
Rh001_037_004+    i_037    tia_h_in_001_004+    5000
Rh001_037_004-    i_037    tia_h_in_001_004-    14736.893704250531
Rh001_038_004+    i_038    tia_h_in_001_004+    13725.297602066792
Rh001_038_004-    i_038    tia_h_in_001_004-    14921.769505094657
Rh001_039_004+    i_039    tia_h_in_001_004+    15000
Rh001_039_004-    i_039    tia_h_in_001_004-    14984.11631830042
Rh001_040_004+    i_040    tia_h_in_001_004+    14802.23828102228
Rh001_040_004-    i_040    tia_h_in_001_004-    15060.834502228581
Rh001_041_004+    i_041    tia_h_in_001_004+    14948.809370880188
Rh001_041_004-    i_041    tia_h_in_001_004-    14889.045398523087
Rh001_042_004+    i_042    tia_h_in_001_004+    14962.590672810868
Rh001_042_004-    i_042    tia_h_in_001_004-    13769.089443781018
Rh001_043_004+    i_043    tia_h_in_001_004+    15135.670976276133
Rh001_043_004-    i_043    tia_h_in_001_004-    13734.47680365261
Rh001_044_004+    i_044    tia_h_in_001_004+    15029.433326921144
Rh001_044_004-    i_044    tia_h_in_001_004-    13644.498789107818
Rh001_045_004+    i_045    tia_h_in_001_004+    14201.947149833066
Rh001_045_004-    i_045    tia_h_in_001_004-    15124.748839552944
Rh001_046_004+    i_046    tia_h_in_001_004+    15101.865249978517
Rh001_046_004-    i_046    tia_h_in_001_004-    14119.195144247966
Rh001_047_004+    i_047    tia_h_in_001_004+    15098.76582316646
Rh001_047_004-    i_047    tia_h_in_001_004-    14569.583970954654
Rh001_048_004+    i_048    tia_h_in_001_004+    15000
Rh001_048_004-    i_048    tia_h_in_001_004-    14138.43954157568
Rh001_049_004+    i_049    tia_h_in_001_004+    14882.635204713866
Rh001_049_004-    i_049    tia_h_in_001_004-    14537.827485426727
Rh001_050_004+    i_050    tia_h_in_001_004+    15012.234980187717
Rh001_050_004-    i_050    tia_h_in_001_004-    13796.05110336512
Rh001_051_004+    i_051    tia_h_in_001_004+    14907.553955588199
Rh001_051_004-    i_051    tia_h_in_001_004-    13967.393572970383
Rh001_052_004+    i_052    tia_h_in_001_004+    14381.280897252194
Rh001_052_004-    i_052    tia_h_in_001_004-    15211.869967472207
Rh001_053_004+    i_053    tia_h_in_001_004+    15058.404935104645
Rh001_053_004-    i_053    tia_h_in_001_004-    14342.772569227853
Rh001_054_004+    i_054    tia_h_in_001_004+    14208.797817605273
Rh001_054_004-    i_054    tia_h_in_001_004-    14804.453456073412
Rh001_055_004+    i_055    tia_h_in_001_004+    15069.497967064954
Rh001_055_004-    i_055    tia_h_in_001_004-    14548.467894116755
Rh001_056_004+    i_056    tia_h_in_001_004+    14863.736510630737
Rh001_056_004-    i_056    tia_h_in_001_004-    13721.280097213652
Rh001_057_004+    i_057    tia_h_in_001_004+    15126.752541509126
Rh001_057_004-    i_057    tia_h_in_001_004-    14532.928927585654
Rh001_058_004+    i_058    tia_h_in_001_004+    15017.391825260913
Rh001_058_004-    i_058    tia_h_in_001_004-    5000
Rh001_059_004+    i_059    tia_h_in_001_004+    15000
Rh001_059_004-    i_059    tia_h_in_001_004-    14383.841587513667
Rh001_060_004+    i_060    tia_h_in_001_004+    14876.95565124784
Rh001_060_004-    i_060    tia_h_in_001_004-    13452.902547313324
Rh001_061_004+    i_061    tia_h_in_001_004+    14232.108908670938
Rh001_061_004-    i_061    tia_h_in_001_004-    15107.303740106165
Rh001_062_004+    i_062    tia_h_in_001_004+    15000
Rh001_062_004-    i_062    tia_h_in_001_004-    13636.717997051861
Rh001_063_004+    i_063    tia_h_in_001_004+    14266.977152392285
Rh001_063_004-    i_063    tia_h_in_001_004-    15159.242222288993
Rh001_064_004+    i_064    tia_h_in_001_004+    14353.472939088877
Rh001_064_004-    i_064    tia_h_in_001_004-    15086.177976118273

* Neuron 5
Rh001_001_005+    i_001    tia_h_in_001_005+    14885.203576538233
Rh001_001_005-    i_001    tia_h_in_001_005-    10975.392450635756
Rh001_002_005+    i_002    tia_h_in_001_005+    14998.637788708851
Rh001_002_005-    i_002    tia_h_in_001_005-    15000
Rh001_003_005+    i_003    tia_h_in_001_005+    14985.29362024385
Rh001_003_005-    i_003    tia_h_in_001_005-    13564.004570059355
Rh001_004_005+    i_004    tia_h_in_001_005+    14798.59007241641
Rh001_004_005-    i_004    tia_h_in_001_005-    12965.230845056947
Rh001_005_005+    i_005    tia_h_in_001_005+    15004.486277384965
Rh001_005_005-    i_005    tia_h_in_001_005-    5000
Rh001_006_005+    i_006    tia_h_in_001_005+    14989.328850581322
Rh001_006_005-    i_006    tia_h_in_001_005-    15203.796330990082
Rh001_007_005+    i_007    tia_h_in_001_005+    15133.284622682339
Rh001_007_005-    i_007    tia_h_in_001_005-    13228.80401919392
Rh001_008_005+    i_008    tia_h_in_001_005+    15053.608592829949
Rh001_008_005-    i_008    tia_h_in_001_005-    14333.781262282817
Rh001_009_005+    i_009    tia_h_in_001_005+    14543.502016434342
Rh001_009_005-    i_009    tia_h_in_001_005-    14798.638017143256
Rh001_010_005+    i_010    tia_h_in_001_005+    10994.800331944494
Rh001_010_005-    i_010    tia_h_in_001_005-    15000
Rh001_011_005+    i_011    tia_h_in_001_005+    5000
Rh001_011_005-    i_011    tia_h_in_001_005-    15152.733734724263
Rh001_012_005+    i_012    tia_h_in_001_005+    14712.458722137855
Rh001_012_005-    i_012    tia_h_in_001_005-    15000
Rh001_013_005+    i_013    tia_h_in_001_005+    13676.935357214626
Rh001_013_005-    i_013    tia_h_in_001_005-    14868.440843639497
Rh001_014_005+    i_014    tia_h_in_001_005+    12413.777870946209
Rh001_014_005-    i_014    tia_h_in_001_005-    15160.573740624026
Rh001_015_005+    i_015    tia_h_in_001_005+    12631.919397471911
Rh001_015_005-    i_015    tia_h_in_001_005-    15000
Rh001_016_005+    i_016    tia_h_in_001_005+    12839.578322282707
Rh001_016_005-    i_016    tia_h_in_001_005-    15010.672802928086
Rh001_017_005+    i_017    tia_h_in_001_005+    15064.64032878056
Rh001_017_005-    i_017    tia_h_in_001_005-    14447.148066882562
Rh001_018_005+    i_018    tia_h_in_001_005+    15092.602371937086
Rh001_018_005-    i_018    tia_h_in_001_005-    14112.265987764304
Rh001_019_005+    i_019    tia_h_in_001_005+    12888.730814442682
Rh001_019_005-    i_019    tia_h_in_001_005-    14954.417246984
Rh001_020_005+    i_020    tia_h_in_001_005+    14990.315032323135
Rh001_020_005-    i_020    tia_h_in_001_005-    15000
Rh001_021_005+    i_021    tia_h_in_001_005+    15156.6297922555
Rh001_021_005-    i_021    tia_h_in_001_005-    13963.568712476637
Rh001_022_005+    i_022    tia_h_in_001_005+    15102.983415378436
Rh001_022_005-    i_022    tia_h_in_001_005-    12623.379831974238
Rh001_023_005+    i_023    tia_h_in_001_005+    15073.778100265412
Rh001_023_005-    i_023    tia_h_in_001_005-    13017.360767167043
Rh001_024_005+    i_024    tia_h_in_001_005+    14337.209169791091
Rh001_024_005-    i_024    tia_h_in_001_005-    14902.342362196068
Rh001_025_005+    i_025    tia_h_in_001_005+    14905.593098384918
Rh001_025_005-    i_025    tia_h_in_001_005-    15059.19654983258
Rh001_026_005+    i_026    tia_h_in_001_005+    14229.722836480483
Rh001_026_005-    i_026    tia_h_in_001_005-    15016.40145881809
Rh001_027_005+    i_027    tia_h_in_001_005+    14160.186903580989
Rh001_027_005-    i_027    tia_h_in_001_005-    14851.243975109848
Rh001_028_005+    i_028    tia_h_in_001_005+    13982.791830463144
Rh001_028_005-    i_028    tia_h_in_001_005-    14881.133850231217
Rh001_029_005+    i_029    tia_h_in_001_005+    15211.633369763063
Rh001_029_005-    i_029    tia_h_in_001_005-    14314.081999492882
Rh001_030_005+    i_030    tia_h_in_001_005+    15100.735883708574
Rh001_030_005-    i_030    tia_h_in_001_005-    13329.751056161407
Rh001_031_005+    i_031    tia_h_in_001_005+    14099.251661900624
Rh001_031_005-    i_031    tia_h_in_001_005-    14956.242628120972
Rh001_032_005+    i_032    tia_h_in_001_005+    5000
Rh001_032_005-    i_032    tia_h_in_001_005-    15000
Rh001_033_005+    i_033    tia_h_in_001_005+    14902.009146899827
Rh001_033_005-    i_033    tia_h_in_001_005-    14123.79152187761
Rh001_034_005+    i_034    tia_h_in_001_005+    14985.587824368415
Rh001_034_005-    i_034    tia_h_in_001_005-    5000
Rh001_035_005+    i_035    tia_h_in_001_005+    14969.15130456166
Rh001_035_005-    i_035    tia_h_in_001_005-    14271.753002565052
Rh001_036_005+    i_036    tia_h_in_001_005+    14864.88429743807
Rh001_036_005-    i_036    tia_h_in_001_005-    15065.538994436169
Rh001_037_005+    i_037    tia_h_in_001_005+    15090.818428224537
Rh001_037_005-    i_037    tia_h_in_001_005-    14896.788746667431
Rh001_038_005+    i_038    tia_h_in_001_005+    14824.140800483101
Rh001_038_005-    i_038    tia_h_in_001_005-    14152.18348966353
Rh001_039_005+    i_039    tia_h_in_001_005+    15103.690147363994
Rh001_039_005-    i_039    tia_h_in_001_005-    13819.08774082371
Rh001_040_005+    i_040    tia_h_in_001_005+    14483.752829432284
Rh001_040_005-    i_040    tia_h_in_001_005-    5000
Rh001_041_005+    i_041    tia_h_in_001_005+    5000
Rh001_041_005-    i_041    tia_h_in_001_005-    15026.778909097333
Rh001_042_005+    i_042    tia_h_in_001_005+    14994.455216708391
Rh001_042_005-    i_042    tia_h_in_001_005-    14457.706774044738
Rh001_043_005+    i_043    tia_h_in_001_005+    15059.692784464884
Rh001_043_005-    i_043    tia_h_in_001_005-    11665.474901517151
Rh001_044_005+    i_044    tia_h_in_001_005+    13525.069802831946
Rh001_044_005-    i_044    tia_h_in_001_005-    15118.127573139145
Rh001_045_005+    i_045    tia_h_in_001_005+    12916.24637473948
Rh001_045_005-    i_045    tia_h_in_001_005-    15075.052935909298
Rh001_046_005+    i_046    tia_h_in_001_005+    5000
Rh001_046_005-    i_046    tia_h_in_001_005-    14559.152879304029
Rh001_047_005+    i_047    tia_h_in_001_005+    14866.47133425165
Rh001_047_005-    i_047    tia_h_in_001_005-    11825.456658312782
Rh001_048_005+    i_048    tia_h_in_001_005+    14934.73363078011
Rh001_048_005-    i_048    tia_h_in_001_005-    13327.61030057908
Rh001_049_005+    i_049    tia_h_in_001_005+    15095.854651932283
Rh001_049_005-    i_049    tia_h_in_001_005-    14522.425757001394
Rh001_050_005+    i_050    tia_h_in_001_005+    14604.385753952429
Rh001_050_005-    i_050    tia_h_in_001_005-    15000
Rh001_051_005+    i_051    tia_h_in_001_005+    13729.011526511636
Rh001_051_005-    i_051    tia_h_in_001_005-    14828.585659329148
Rh001_052_005+    i_052    tia_h_in_001_005+    14862.244187074768
Rh001_052_005-    i_052    tia_h_in_001_005-    13411.512176493487
Rh001_053_005+    i_053    tia_h_in_001_005+    15000
Rh001_053_005-    i_053    tia_h_in_001_005-    15351.927856125201
Rh001_054_005+    i_054    tia_h_in_001_005+    12936.862814488406
Rh001_054_005-    i_054    tia_h_in_001_005-    15132.036929496864
Rh001_055_005+    i_055    tia_h_in_001_005+    12639.136765403631
Rh001_055_005-    i_055    tia_h_in_001_005-    15139.473583272844
Rh001_056_005+    i_056    tia_h_in_001_005+    15034.291226959282
Rh001_056_005-    i_056    tia_h_in_001_005-    13593.455642854278
Rh001_057_005+    i_057    tia_h_in_001_005+    13700.10185666359
Rh001_057_005-    i_057    tia_h_in_001_005-    15017.207620153014
Rh001_058_005+    i_058    tia_h_in_001_005+    15000
Rh001_058_005-    i_058    tia_h_in_001_005-    5000
Rh001_059_005+    i_059    tia_h_in_001_005+    13873.555006533861
Rh001_059_005-    i_059    tia_h_in_001_005-    15082.531732684194
Rh001_060_005+    i_060    tia_h_in_001_005+    14727.79464200269
Rh001_060_005-    i_060    tia_h_in_001_005-    15164.068486359178
Rh001_061_005+    i_061    tia_h_in_001_005+    14999.64463363475
Rh001_061_005-    i_061    tia_h_in_001_005-    13751.889001298261
Rh001_062_005+    i_062    tia_h_in_001_005+    14027.681146529183
Rh001_062_005-    i_062    tia_h_in_001_005-    15123.182952405392
Rh001_063_005+    i_063    tia_h_in_001_005+    11693.927218842216
Rh001_063_005-    i_063    tia_h_in_001_005-    14883.406287788348
Rh001_064_005+    i_064    tia_h_in_001_005+    15018.782645577994
Rh001_064_005-    i_064    tia_h_in_001_005-    12256.716695632846

* Neuron 6
Rh001_001_006+    i_001    tia_h_in_001_006+    14992.106092693113
Rh001_001_006-    i_001    tia_h_in_001_006-    14100.356953691593
Rh001_002_006+    i_002    tia_h_in_001_006+    14864.020574073655
Rh001_002_006-    i_002    tia_h_in_001_006-    13676.97794827337
Rh001_003_006+    i_003    tia_h_in_001_006+    14970.352127733098
Rh001_003_006-    i_003    tia_h_in_001_006-    13834.583989507935
Rh001_004_006+    i_004    tia_h_in_001_006+    15034.451109034613
Rh001_004_006-    i_004    tia_h_in_001_006-    13601.996382191242
Rh001_005_006+    i_005    tia_h_in_001_006+    14871.047709450593
Rh001_005_006-    i_005    tia_h_in_001_006-    13668.938399913222
Rh001_006_006+    i_006    tia_h_in_001_006+    15212.438661916505
Rh001_006_006-    i_006    tia_h_in_001_006-    14382.541457787811
Rh001_007_006+    i_007    tia_h_in_001_006+    15000
Rh001_007_006-    i_007    tia_h_in_001_006-    15052.445981373541
Rh001_008_006+    i_008    tia_h_in_001_006+    5000
Rh001_008_006-    i_008    tia_h_in_001_006-    15022.52101915787
Rh001_009_006+    i_009    tia_h_in_001_006+    15034.467484580291
Rh001_009_006-    i_009    tia_h_in_001_006-    13879.387875248918
Rh001_010_006+    i_010    tia_h_in_001_006+    14991.350202999447
Rh001_010_006-    i_010    tia_h_in_001_006-    13662.09597213927
Rh001_011_006+    i_011    tia_h_in_001_006+    14401.483285530188
Rh001_011_006-    i_011    tia_h_in_001_006-    14872.412681847345
Rh001_012_006+    i_012    tia_h_in_001_006+    15253.463161634103
Rh001_012_006-    i_012    tia_h_in_001_006-    13619.707063702637
Rh001_013_006+    i_013    tia_h_in_001_006+    14976.252479778952
Rh001_013_006-    i_013    tia_h_in_001_006-    14531.737146833073
Rh001_014_006+    i_014    tia_h_in_001_006+    14367.781228089014
Rh001_014_006-    i_014    tia_h_in_001_006-    5000
Rh001_015_006+    i_015    tia_h_in_001_006+    15080.300530499684
Rh001_015_006-    i_015    tia_h_in_001_006-    14137.97167115076
Rh001_016_006+    i_016    tia_h_in_001_006+    14894.766038782187
Rh001_016_006-    i_016    tia_h_in_001_006-    14720.867154197995
Rh001_017_006+    i_017    tia_h_in_001_006+    14916.283852159295
Rh001_017_006-    i_017    tia_h_in_001_006-    14878.578904496717
Rh001_018_006+    i_018    tia_h_in_001_006+    15055.460335094127
Rh001_018_006-    i_018    tia_h_in_001_006-    14551.361302615112
Rh001_019_006+    i_019    tia_h_in_001_006+    15291.4746805687
Rh001_019_006-    i_019    tia_h_in_001_006-    14059.591933232408
Rh001_020_006+    i_020    tia_h_in_001_006+    14812.44832427093
Rh001_020_006-    i_020    tia_h_in_001_006-    13457.737109909278
Rh001_021_006+    i_021    tia_h_in_001_006+    14860.922406587893
Rh001_021_006-    i_021    tia_h_in_001_006-    13804.815604911299
Rh001_022_006+    i_022    tia_h_in_001_006+    15033.766129077418
Rh001_022_006-    i_022    tia_h_in_001_006-    14116.805082631403
Rh001_023_006+    i_023    tia_h_in_001_006+    13695.25789048949
Rh001_023_006-    i_023    tia_h_in_001_006-    15090.118241306865
Rh001_024_006+    i_024    tia_h_in_001_006+    15192.52713162286
Rh001_024_006-    i_024    tia_h_in_001_006-    14168.31747227878
Rh001_025_006+    i_025    tia_h_in_001_006+    15129.598934945241
Rh001_025_006-    i_025    tia_h_in_001_006-    14049.73143113946
Rh001_026_006+    i_026    tia_h_in_001_006+    14524.139554529973
Rh001_026_006-    i_026    tia_h_in_001_006-    15003.377777822883
Rh001_027_006+    i_027    tia_h_in_001_006+    14722.464299707228
Rh001_027_006-    i_027    tia_h_in_001_006-    14968.204706455323
Rh001_028_006+    i_028    tia_h_in_001_006+    14300.547788852662
Rh001_028_006-    i_028    tia_h_in_001_006-    14951.325824835405
Rh001_029_006+    i_029    tia_h_in_001_006+    13840.312957322249
Rh001_029_006-    i_029    tia_h_in_001_006-    14907.347942588254
Rh001_030_006+    i_030    tia_h_in_001_006+    13958.91213929624
Rh001_030_006-    i_030    tia_h_in_001_006-    14987.028401410107
Rh001_031_006+    i_031    tia_h_in_001_006+    14959.387708141645
Rh001_031_006-    i_031    tia_h_in_001_006-    13256.340303606969
Rh001_032_006+    i_032    tia_h_in_001_006+    14931.464302109427
Rh001_032_006-    i_032    tia_h_in_001_006-    14992.343384737736
Rh001_033_006+    i_033    tia_h_in_001_006+    13949.492625346922
Rh001_033_006-    i_033    tia_h_in_001_006-    15122.715093564853
Rh001_034_006+    i_034    tia_h_in_001_006+    15122.074480025303
Rh001_034_006-    i_034    tia_h_in_001_006-    14501.414085492603
Rh001_035_006+    i_035    tia_h_in_001_006+    15049.618863715064
Rh001_035_006-    i_035    tia_h_in_001_006-    13939.686469253262
Rh001_036_006+    i_036    tia_h_in_001_006+    13487.679741456219
Rh001_036_006-    i_036    tia_h_in_001_006-    15120.322363990095
Rh001_037_006+    i_037    tia_h_in_001_006+    15012.33735778924
Rh001_037_006-    i_037    tia_h_in_001_006-    14138.728646098656
Rh001_038_006+    i_038    tia_h_in_001_006+    14766.64705611708
Rh001_038_006-    i_038    tia_h_in_001_006-    14092.903107450631
Rh001_039_006+    i_039    tia_h_in_001_006+    15122.759077177265
Rh001_039_006-    i_039    tia_h_in_001_006-    13637.899385820123
Rh001_040_006+    i_040    tia_h_in_001_006+    15030.690673123992
Rh001_040_006-    i_040    tia_h_in_001_006-    15093.462472555791
Rh001_041_006+    i_041    tia_h_in_001_006+    14553.65363565243
Rh001_041_006-    i_041    tia_h_in_001_006-    15137.219318524627
Rh001_042_006+    i_042    tia_h_in_001_006+    14824.239923685464
Rh001_042_006-    i_042    tia_h_in_001_006-    14917.275119413649
Rh001_043_006+    i_043    tia_h_in_001_006+    15000
Rh001_043_006-    i_043    tia_h_in_001_006-    15044.425419375386
Rh001_044_006+    i_044    tia_h_in_001_006+    15090.267848405587
Rh001_044_006-    i_044    tia_h_in_001_006-    13828.406165103223
Rh001_045_006+    i_045    tia_h_in_001_006+    15146.044221374985
Rh001_045_006-    i_045    tia_h_in_001_006-    13588.459279517407
Rh001_046_006+    i_046    tia_h_in_001_006+    14954.851685394191
Rh001_046_006-    i_046    tia_h_in_001_006-    14899.6555963466
Rh001_047_006+    i_047    tia_h_in_001_006+    13730.195797577762
Rh001_047_006-    i_047    tia_h_in_001_006-    5000
Rh001_048_006+    i_048    tia_h_in_001_006+    15000
Rh001_048_006-    i_048    tia_h_in_001_006-    14960.80391939456
Rh001_049_006+    i_049    tia_h_in_001_006+    15250.424933073544
Rh001_049_006-    i_049    tia_h_in_001_006-    14020.401167004426
Rh001_050_006+    i_050    tia_h_in_001_006+    14774.232757227983
Rh001_050_006-    i_050    tia_h_in_001_006-    15039.599706835985
Rh001_051_006+    i_051    tia_h_in_001_006+    15033.732462411792
Rh001_051_006-    i_051    tia_h_in_001_006-    13981.02689700276
Rh001_052_006+    i_052    tia_h_in_001_006+    15013.031235233475
Rh001_052_006-    i_052    tia_h_in_001_006-    14222.42263034504
Rh001_053_006+    i_053    tia_h_in_001_006+    14938.88845766233
Rh001_053_006-    i_053    tia_h_in_001_006-    14986.9938438236
Rh001_054_006+    i_054    tia_h_in_001_006+    14447.143476359568
Rh001_054_006-    i_054    tia_h_in_001_006-    14933.9565462599
Rh001_055_006+    i_055    tia_h_in_001_006+    13747.978609423437
Rh001_055_006-    i_055    tia_h_in_001_006-    14862.403435095974
Rh001_056_006+    i_056    tia_h_in_001_006+    15005.800640692958
Rh001_056_006-    i_056    tia_h_in_001_006-    13639.149682563937
Rh001_057_006+    i_057    tia_h_in_001_006+    14057.880376325656
Rh001_057_006-    i_057    tia_h_in_001_006-    15099.441663705133
Rh001_058_006+    i_058    tia_h_in_001_006+    15014.90483034529
Rh001_058_006-    i_058    tia_h_in_001_006-    5000
Rh001_059_006+    i_059    tia_h_in_001_006+    15000
Rh001_059_006-    i_059    tia_h_in_001_006-    14973.995109315141
Rh001_060_006+    i_060    tia_h_in_001_006+    13920.418239792318
Rh001_060_006-    i_060    tia_h_in_001_006-    14827.80321537867
Rh001_061_006+    i_061    tia_h_in_001_006+    14973.608531287764
Rh001_061_006-    i_061    tia_h_in_001_006-    15041.660251631649
Rh001_062_006+    i_062    tia_h_in_001_006+    13924.470574825787
Rh001_062_006-    i_062    tia_h_in_001_006-    15245.610852263735
Rh001_063_006+    i_063    tia_h_in_001_006+    15121.976659105429
Rh001_063_006-    i_063    tia_h_in_001_006-    13563.99412925854
Rh001_064_006+    i_064    tia_h_in_001_006+    14883.237830249876
Rh001_064_006-    i_064    tia_h_in_001_006-    15000

* Neuron 7
Rh001_001_007+    i_001    tia_h_in_001_007+    13713.67563164278
Rh001_001_007-    i_001    tia_h_in_001_007-    15080.312684469269
Rh001_002_007+    i_002    tia_h_in_001_007+    5000
Rh001_002_007-    i_002    tia_h_in_001_007-    14621.736039892827
Rh001_003_007+    i_003    tia_h_in_001_007+    14799.519908835633
Rh001_003_007-    i_003    tia_h_in_001_007-    14437.573179739198
Rh001_004_007+    i_004    tia_h_in_001_007+    13070.92738969988
Rh001_004_007-    i_004    tia_h_in_001_007-    14885.5919044148
Rh001_005_007+    i_005    tia_h_in_001_007+    14191.072212505826
Rh001_005_007-    i_005    tia_h_in_001_007-    15037.474045116598
Rh001_006_007+    i_006    tia_h_in_001_007+    14433.030157122732
Rh001_006_007-    i_006    tia_h_in_001_007-    15017.857223701392
Rh001_007_007+    i_007    tia_h_in_001_007+    13654.906680016675
Rh001_007_007-    i_007    tia_h_in_001_007-    14991.451053542163
Rh001_008_007+    i_008    tia_h_in_001_007+    13941.900007917715
Rh001_008_007-    i_008    tia_h_in_001_007-    15025.659752664975
Rh001_009_007+    i_009    tia_h_in_001_007+    14992.150070493686
Rh001_009_007-    i_009    tia_h_in_001_007-    11769.991816557304
Rh001_010_007+    i_010    tia_h_in_001_007+    14989.630416326618
Rh001_010_007-    i_010    tia_h_in_001_007-    13371.57398229572
Rh001_011_007+    i_011    tia_h_in_001_007+    12991.018322995957
Rh001_011_007-    i_011    tia_h_in_001_007-    15184.276101985393
Rh001_012_007+    i_012    tia_h_in_001_007+    15000
Rh001_012_007-    i_012    tia_h_in_001_007-    14964.612648441278
Rh001_013_007+    i_013    tia_h_in_001_007+    15064.348474868228
Rh001_013_007-    i_013    tia_h_in_001_007-    15075.862040754344
Rh001_014_007+    i_014    tia_h_in_001_007+    12895.174107738323
Rh001_014_007-    i_014    tia_h_in_001_007-    15099.750353077572
Rh001_015_007+    i_015    tia_h_in_001_007+    14216.526281346649
Rh001_015_007-    i_015    tia_h_in_001_007-    15000
Rh001_016_007+    i_016    tia_h_in_001_007+    12903.008894461054
Rh001_016_007-    i_016    tia_h_in_001_007-    14942.532803441101
Rh001_017_007+    i_017    tia_h_in_001_007+    15002.719504581522
Rh001_017_007-    i_017    tia_h_in_001_007-    13314.438632955858
Rh001_018_007+    i_018    tia_h_in_001_007+    15000
Rh001_018_007-    i_018    tia_h_in_001_007-    13403.089293298535
Rh001_019_007+    i_019    tia_h_in_001_007+    5000
Rh001_019_007-    i_019    tia_h_in_001_007-    12507.2871923354
Rh001_020_007+    i_020    tia_h_in_001_007+    15063.880160486091
Rh001_020_007-    i_020    tia_h_in_001_007-    14489.62908135321
Rh001_021_007+    i_021    tia_h_in_001_007+    14663.354608268959
Rh001_021_007-    i_021    tia_h_in_001_007-    14220.43151353909
Rh001_022_007+    i_022    tia_h_in_001_007+    14951.90022494095
Rh001_022_007-    i_022    tia_h_in_001_007-    12866.626377887082
Rh001_023_007+    i_023    tia_h_in_001_007+    14905.437198547344
Rh001_023_007-    i_023    tia_h_in_001_007-    15000
Rh001_024_007+    i_024    tia_h_in_001_007+    14873.348283419009
Rh001_024_007-    i_024    tia_h_in_001_007-    15055.36183756545
Rh001_025_007+    i_025    tia_h_in_001_007+    13955.954822391246
Rh001_025_007-    i_025    tia_h_in_001_007-    5000
Rh001_026_007+    i_026    tia_h_in_001_007+    12554.609663565037
Rh001_026_007-    i_026    tia_h_in_001_007-    14959.306530049473
Rh001_027_007+    i_027    tia_h_in_001_007+    14941.349469173505
Rh001_027_007-    i_027    tia_h_in_001_007-    15022.151342481384
Rh001_028_007+    i_028    tia_h_in_001_007+    14841.305815787158
Rh001_028_007-    i_028    tia_h_in_001_007-    14070.121237684418
Rh001_029_007+    i_029    tia_h_in_001_007+    14920.981763191992
Rh001_029_007-    i_029    tia_h_in_001_007-    13396.577820895907
Rh001_030_007+    i_030    tia_h_in_001_007+    14774.232733911169
Rh001_030_007-    i_030    tia_h_in_001_007-    14704.834014671582
Rh001_031_007+    i_031    tia_h_in_001_007+    14959.203006101623
Rh001_031_007-    i_031    tia_h_in_001_007-    14176.283029935159
Rh001_032_007+    i_032    tia_h_in_001_007+    15093.488333060703
Rh001_032_007-    i_032    tia_h_in_001_007-    14199.694466733084
Rh001_033_007+    i_033    tia_h_in_001_007+    14795.208575626946
Rh001_033_007-    i_033    tia_h_in_001_007-    15174.663706906638
Rh001_034_007+    i_034    tia_h_in_001_007+    13357.692029502172
Rh001_034_007-    i_034    tia_h_in_001_007-    15059.877834608244
Rh001_035_007+    i_035    tia_h_in_001_007+    15000
Rh001_035_007-    i_035    tia_h_in_001_007-    12080.950555699437
Rh001_036_007+    i_036    tia_h_in_001_007+    5000
Rh001_036_007-    i_036    tia_h_in_001_007-    14709.483919482427
Rh001_037_007+    i_037    tia_h_in_001_007+    13989.629182067987
Rh001_037_007-    i_037    tia_h_in_001_007-    14962.27841994812
Rh001_038_007+    i_038    tia_h_in_001_007+    14893.02084310729
Rh001_038_007-    i_038    tia_h_in_001_007-    13243.220037205974
Rh001_039_007+    i_039    tia_h_in_001_007+    13907.419903260867
Rh001_039_007-    i_039    tia_h_in_001_007-    15212.544215742495
Rh001_040_007+    i_040    tia_h_in_001_007+    15046.71849783262
Rh001_040_007-    i_040    tia_h_in_001_007-    13570.84677019603
Rh001_041_007+    i_041    tia_h_in_001_007+    5000
Rh001_041_007-    i_041    tia_h_in_001_007-    15177.887915792762
Rh001_042_007+    i_042    tia_h_in_001_007+    13801.92360605778
Rh001_042_007-    i_042    tia_h_in_001_007-    15195.579186248446
Rh001_043_007+    i_043    tia_h_in_001_007+    15121.792850464786
Rh001_043_007-    i_043    tia_h_in_001_007-    5000
Rh001_044_007+    i_044    tia_h_in_001_007+    14469.255889209555
Rh001_044_007-    i_044    tia_h_in_001_007-    15020.567317534744
Rh001_045_007+    i_045    tia_h_in_001_007+    15100.635376788356
Rh001_045_007-    i_045    tia_h_in_001_007-    12808.013853035667
Rh001_046_007+    i_046    tia_h_in_001_007+    14739.363619847203
Rh001_046_007-    i_046    tia_h_in_001_007-    5000
Rh001_047_007+    i_047    tia_h_in_001_007+    13431.54111106866
Rh001_047_007-    i_047    tia_h_in_001_007-    5000
Rh001_048_007+    i_048    tia_h_in_001_007+    14586.403327208804
Rh001_048_007-    i_048    tia_h_in_001_007-    15029.069227779833
Rh001_049_007+    i_049    tia_h_in_001_007+    5000
Rh001_049_007-    i_049    tia_h_in_001_007-    14847.204413882113
Rh001_050_007+    i_050    tia_h_in_001_007+    14429.147078653925
Rh001_050_007-    i_050    tia_h_in_001_007-    14958.464233866687
Rh001_051_007+    i_051    tia_h_in_001_007+    11979.513113932342
Rh001_051_007-    i_051    tia_h_in_001_007-    14927.937124631659
Rh001_052_007+    i_052    tia_h_in_001_007+    15000
Rh001_052_007-    i_052    tia_h_in_001_007-    14892.87274252013
Rh001_053_007+    i_053    tia_h_in_001_007+    12635.636049651957
Rh001_053_007-    i_053    tia_h_in_001_007-    14968.62543295425
Rh001_054_007+    i_054    tia_h_in_001_007+    11141.626730243974
Rh001_054_007-    i_054    tia_h_in_001_007-    15077.79963274839
Rh001_055_007+    i_055    tia_h_in_001_007+    12323.141051985089
Rh001_055_007-    i_055    tia_h_in_001_007-    15138.04261265524
Rh001_056_007+    i_056    tia_h_in_001_007+    13448.633694311244
Rh001_056_007-    i_056    tia_h_in_001_007-    15212.7504491324
Rh001_057_007+    i_057    tia_h_in_001_007+    13750.541013607211
Rh001_057_007-    i_057    tia_h_in_001_007-    15000
Rh001_058_007+    i_058    tia_h_in_001_007+    15127.396059444865
Rh001_058_007-    i_058    tia_h_in_001_007-    14324.212574661837
Rh001_059_007+    i_059    tia_h_in_001_007+    14916.252010341386
Rh001_059_007-    i_059    tia_h_in_001_007-    12936.416377635749
Rh001_060_007+    i_060    tia_h_in_001_007+    14935.896445357414
Rh001_060_007-    i_060    tia_h_in_001_007-    15000
Rh001_061_007+    i_061    tia_h_in_001_007+    13917.449493000551
Rh001_061_007-    i_061    tia_h_in_001_007-    14913.285139431302
Rh001_062_007+    i_062    tia_h_in_001_007+    15000
Rh001_062_007-    i_062    tia_h_in_001_007-    10772.963321601062
Rh001_063_007+    i_063    tia_h_in_001_007+    15000
Rh001_063_007-    i_063    tia_h_in_001_007-    10034.585566587482
Rh001_064_007+    i_064    tia_h_in_001_007+    14819.025480209604
Rh001_064_007-    i_064    tia_h_in_001_007-    5000

* Neuron 8
Rh001_001_008+    i_001    tia_h_in_001_008+    14858.267968032045
Rh001_001_008-    i_001    tia_h_in_001_008-    12756.309502918002
Rh001_002_008+    i_002    tia_h_in_001_008+    13249.6971204251
Rh001_002_008-    i_002    tia_h_in_001_008-    14725.520017133851
Rh001_003_008+    i_003    tia_h_in_001_008+    14949.61143628452
Rh001_003_008-    i_003    tia_h_in_001_008-    13794.605796630702
Rh001_004_008+    i_004    tia_h_in_001_008+    15000
Rh001_004_008-    i_004    tia_h_in_001_008-    14398.339642487259
Rh001_005_008+    i_005    tia_h_in_001_008+    14843.974765837931
Rh001_005_008-    i_005    tia_h_in_001_008-    15002.79223261231
Rh001_006_008+    i_006    tia_h_in_001_008+    13249.636797489606
Rh001_006_008-    i_006    tia_h_in_001_008-    14995.212382785177
Rh001_007_008+    i_007    tia_h_in_001_008+    14402.30652839994
Rh001_007_008-    i_007    tia_h_in_001_008-    15118.555556772239
Rh001_008_008+    i_008    tia_h_in_001_008+    12115.953310011739
Rh001_008_008-    i_008    tia_h_in_001_008-    15054.957370951272
Rh001_009_008+    i_009    tia_h_in_001_008+    14304.381527777388
Rh001_009_008-    i_009    tia_h_in_001_008-    14790.500891439879
Rh001_010_008+    i_010    tia_h_in_001_008+    14541.119420741072
Rh001_010_008-    i_010    tia_h_in_001_008-    15083.436694528751
Rh001_011_008+    i_011    tia_h_in_001_008+    13209.28961922685
Rh001_011_008-    i_011    tia_h_in_001_008-    15107.479956072355
Rh001_012_008+    i_012    tia_h_in_001_008+    14968.363008859347
Rh001_012_008-    i_012    tia_h_in_001_008-    12281.83521515919
Rh001_013_008+    i_013    tia_h_in_001_008+    14949.397936661404
Rh001_013_008-    i_013    tia_h_in_001_008-    14442.332324582097
Rh001_014_008+    i_014    tia_h_in_001_008+    14874.986659525226
Rh001_014_008-    i_014    tia_h_in_001_008-    13493.278709397733
Rh001_015_008+    i_015    tia_h_in_001_008+    15011.71683233584
Rh001_015_008-    i_015    tia_h_in_001_008-    15000
Rh001_016_008+    i_016    tia_h_in_001_008+    15155.722961554482
Rh001_016_008-    i_016    tia_h_in_001_008-    14522.289063491913
Rh001_017_008+    i_017    tia_h_in_001_008+    12237.65384711669
Rh001_017_008-    i_017    tia_h_in_001_008-    14876.5514997407
Rh001_018_008+    i_018    tia_h_in_001_008+    13701.202590979214
Rh001_018_008-    i_018    tia_h_in_001_008-    14969.774340689892
Rh001_019_008+    i_019    tia_h_in_001_008+    12274.832644802573
Rh001_019_008-    i_019    tia_h_in_001_008-    14972.210852178358
Rh001_020_008+    i_020    tia_h_in_001_008+    12113.961325151813
Rh001_020_008-    i_020    tia_h_in_001_008-    14953.908598780898
Rh001_021_008+    i_021    tia_h_in_001_008+    13782.585200100852
Rh001_021_008-    i_021    tia_h_in_001_008-    15129.628931789084
Rh001_022_008+    i_022    tia_h_in_001_008+    15203.848882896937
Rh001_022_008-    i_022    tia_h_in_001_008-    13219.53083702607
Rh001_023_008+    i_023    tia_h_in_001_008+    14646.363079470457
Rh001_023_008-    i_023    tia_h_in_001_008-    15000
Rh001_024_008+    i_024    tia_h_in_001_008+    14947.218803690013
Rh001_024_008-    i_024    tia_h_in_001_008-    11878.842504744918
Rh001_025_008+    i_025    tia_h_in_001_008+    14777.175586893021
Rh001_025_008-    i_025    tia_h_in_001_008-    14916.64657811073
Rh001_026_008+    i_026    tia_h_in_001_008+    15054.018533398516
Rh001_026_008-    i_026    tia_h_in_001_008-    13651.090064336857
Rh001_027_008+    i_027    tia_h_in_001_008+    14302.130396538278
Rh001_027_008-    i_027    tia_h_in_001_008-    14999.895851612548
Rh001_028_008+    i_028    tia_h_in_001_008+    12692.151895149413
Rh001_028_008-    i_028    tia_h_in_001_008-    15072.020228007326
Rh001_029_008+    i_029    tia_h_in_001_008+    15156.254190263302
Rh001_029_008-    i_029    tia_h_in_001_008-    14504.98383293334
Rh001_030_008+    i_030    tia_h_in_001_008+    14923.088997900606
Rh001_030_008-    i_030    tia_h_in_001_008-    15116.222208154539
Rh001_031_008+    i_031    tia_h_in_001_008+    14848.774957025738
Rh001_031_008-    i_031    tia_h_in_001_008-    15000
Rh001_032_008+    i_032    tia_h_in_001_008+    14848.342073298669
Rh001_032_008-    i_032    tia_h_in_001_008-    14622.986503008035
Rh001_033_008+    i_033    tia_h_in_001_008+    15079.543291032267
Rh001_033_008-    i_033    tia_h_in_001_008-    13863.573260989675
Rh001_034_008+    i_034    tia_h_in_001_008+    14037.154232114326
Rh001_034_008-    i_034    tia_h_in_001_008-    15000
Rh001_035_008+    i_035    tia_h_in_001_008+    14551.977798782918
Rh001_035_008-    i_035    tia_h_in_001_008-    15138.536530599393
Rh001_036_008+    i_036    tia_h_in_001_008+    14893.69754171478
Rh001_036_008-    i_036    tia_h_in_001_008-    12357.794950102
Rh001_037_008+    i_037    tia_h_in_001_008+    13679.553323473634
Rh001_037_008-    i_037    tia_h_in_001_008-    15116.47386538227
Rh001_038_008+    i_038    tia_h_in_001_008+    13400.350271178699
Rh001_038_008-    i_038    tia_h_in_001_008-    15094.241806233955
Rh001_039_008+    i_039    tia_h_in_001_008+    14868.979056870738
Rh001_039_008-    i_039    tia_h_in_001_008-    14902.076505781673
Rh001_040_008+    i_040    tia_h_in_001_008+    13303.629391223863
Rh001_040_008-    i_040    tia_h_in_001_008-    15002.09393861688
Rh001_041_008+    i_041    tia_h_in_001_008+    15160.071672438466
Rh001_041_008-    i_041    tia_h_in_001_008-    13593.694319167722
Rh001_042_008+    i_042    tia_h_in_001_008+    15066.923292479458
Rh001_042_008-    i_042    tia_h_in_001_008-    12090.166940283465
Rh001_043_008+    i_043    tia_h_in_001_008+    14991.176491841208
Rh001_043_008-    i_043    tia_h_in_001_008-    13289.718756307502
Rh001_044_008+    i_044    tia_h_in_001_008+    15236.018186094403
Rh001_044_008-    i_044    tia_h_in_001_008-    13111.590315468029
Rh001_045_008+    i_045    tia_h_in_001_008+    14373.05073355177
Rh001_045_008-    i_045    tia_h_in_001_008-    15167.821884138744
Rh001_046_008+    i_046    tia_h_in_001_008+    12335.137222446503
Rh001_046_008-    i_046    tia_h_in_001_008-    14890.675155098588
Rh001_047_008+    i_047    tia_h_in_001_008+    13695.167659295928
Rh001_047_008-    i_047    tia_h_in_001_008-    15070.84317219293
Rh001_048_008+    i_048    tia_h_in_001_008+    11213.778467216904
Rh001_048_008-    i_048    tia_h_in_001_008-    14874.751806756865
Rh001_049_008+    i_049    tia_h_in_001_008+    15006.11522447895
Rh001_049_008-    i_049    tia_h_in_001_008-    14132.905566673477
Rh001_050_008+    i_050    tia_h_in_001_008+    14214.986729570419
Rh001_050_008-    i_050    tia_h_in_001_008-    14932.30954876207
Rh001_051_008+    i_051    tia_h_in_001_008+    14660.2121686253
Rh001_051_008-    i_051    tia_h_in_001_008-    15214.646449064514
Rh001_052_008+    i_052    tia_h_in_001_008+    13397.026098473694
Rh001_052_008-    i_052    tia_h_in_001_008-    14905.919529879366
Rh001_053_008+    i_053    tia_h_in_001_008+    5000
Rh001_053_008-    i_053    tia_h_in_001_008-    14867.654075714003
Rh001_054_008+    i_054    tia_h_in_001_008+    11962.730321505864
Rh001_054_008-    i_054    tia_h_in_001_008-    15019.497252151676
Rh001_055_008+    i_055    tia_h_in_001_008+    11584.46869603379
Rh001_055_008-    i_055    tia_h_in_001_008-    15282.010974802923
Rh001_056_008+    i_056    tia_h_in_001_008+    13942.985087622728
Rh001_056_008-    i_056    tia_h_in_001_008-    14805.98044793599
Rh001_057_008+    i_057    tia_h_in_001_008+    15183.131635709065
Rh001_057_008-    i_057    tia_h_in_001_008-    15027.125259306353
Rh001_058_008+    i_058    tia_h_in_001_008+    14993.008068064506
Rh001_058_008-    i_058    tia_h_in_001_008-    14615.83542866354
Rh001_059_008+    i_059    tia_h_in_001_008+    14471.19673058446
Rh001_059_008-    i_059    tia_h_in_001_008-    14889.310747958652
Rh001_060_008+    i_060    tia_h_in_001_008+    14912.028273639362
Rh001_060_008-    i_060    tia_h_in_001_008-    10764.704961771207
Rh001_061_008+    i_061    tia_h_in_001_008+    15037.602851104977
Rh001_061_008-    i_061    tia_h_in_001_008-    12524.7050064279
Rh001_062_008+    i_062    tia_h_in_001_008+    15000
Rh001_062_008-    i_062    tia_h_in_001_008-    11464.75099290297
Rh001_063_008+    i_063    tia_h_in_001_008+    15153.171008855794
Rh001_063_008-    i_063    tia_h_in_001_008-    9459.432258323539
Rh001_064_008+    i_064    tia_h_in_001_008+    15100.310875989899
Rh001_064_008-    i_064    tia_h_in_001_008-    9673.642588848796

* Neuron 9
Rh001_001_009+    i_001    tia_h_in_001_009+    13809.878215865809
Rh001_001_009-    i_001    tia_h_in_001_009-    15000
Rh001_002_009+    i_002    tia_h_in_001_009+    14873.579570127196
Rh001_002_009-    i_002    tia_h_in_001_009-    12621.388419096513
Rh001_003_009+    i_003    tia_h_in_001_009+    15068.523006794632
Rh001_003_009-    i_003    tia_h_in_001_009-    14486.904338348824
Rh001_004_009+    i_004    tia_h_in_001_009+    14428.993891806746
Rh001_004_009-    i_004    tia_h_in_001_009-    15052.599320017765
Rh001_005_009+    i_005    tia_h_in_001_009+    14786.41363374334
Rh001_005_009-    i_005    tia_h_in_001_009-    14944.814796713528
Rh001_006_009+    i_006    tia_h_in_001_009+    13988.457851909743
Rh001_006_009-    i_006    tia_h_in_001_009-    14890.770090335782
Rh001_007_009+    i_007    tia_h_in_001_009+    15000
Rh001_007_009-    i_007    tia_h_in_001_009-    14996.46724398301
Rh001_008_009+    i_008    tia_h_in_001_009+    5000
Rh001_008_009-    i_008    tia_h_in_001_009-    15039.130957297926
Rh001_009_009+    i_009    tia_h_in_001_009+    5000
Rh001_009_009-    i_009    tia_h_in_001_009-    15025.079773261741
Rh001_010_009+    i_010    tia_h_in_001_009+    14847.189265002628
Rh001_010_009-    i_010    tia_h_in_001_009-    13925.076340429801
Rh001_011_009+    i_011    tia_h_in_001_009+    14471.977384094325
Rh001_011_009-    i_011    tia_h_in_001_009-    14903.263775992158
Rh001_012_009+    i_012    tia_h_in_001_009+    13417.038816451179
Rh001_012_009-    i_012    tia_h_in_001_009-    15071.289883395768
Rh001_013_009+    i_013    tia_h_in_001_009+    15035.715027892713
Rh001_013_009-    i_013    tia_h_in_001_009-    13893.055060186081
Rh001_014_009+    i_014    tia_h_in_001_009+    14846.14742052575
Rh001_014_009-    i_014    tia_h_in_001_009-    15000
Rh001_015_009+    i_015    tia_h_in_001_009+    15109.85773109342
Rh001_015_009-    i_015    tia_h_in_001_009-    13984.5477465881
Rh001_016_009+    i_016    tia_h_in_001_009+    15027.349928807733
Rh001_016_009-    i_016    tia_h_in_001_009-    11787.374144530357
Rh001_017_009+    i_017    tia_h_in_001_009+    5000
Rh001_017_009-    i_017    tia_h_in_001_009-    15000
Rh001_018_009+    i_018    tia_h_in_001_009+    11731.702067736744
Rh001_018_009-    i_018    tia_h_in_001_009-    15038.796273093098
Rh001_019_009+    i_019    tia_h_in_001_009+    14520.066853603563
Rh001_019_009-    i_019    tia_h_in_001_009-    14979.325763673
Rh001_020_009+    i_020    tia_h_in_001_009+    14964.30927783267
Rh001_020_009-    i_020    tia_h_in_001_009-    14440.657346405136
Rh001_021_009+    i_021    tia_h_in_001_009+    15029.800164690254
Rh001_021_009-    i_021    tia_h_in_001_009-    13318.048413979375
Rh001_022_009+    i_022    tia_h_in_001_009+    15020.98464716291
Rh001_022_009-    i_022    tia_h_in_001_009-    5000
Rh001_023_009+    i_023    tia_h_in_001_009+    14992.934472452005
Rh001_023_009-    i_023    tia_h_in_001_009-    14946.511679872248
Rh001_024_009+    i_024    tia_h_in_001_009+    13609.576909808815
Rh001_024_009-    i_024    tia_h_in_001_009-    14940.756514997769
Rh001_025_009+    i_025    tia_h_in_001_009+    15033.638463851556
Rh001_025_009-    i_025    tia_h_in_001_009-    11468.936589241228
Rh001_026_009+    i_026    tia_h_in_001_009+    14856.261688747965
Rh001_026_009-    i_026    tia_h_in_001_009-    14802.888708622939
Rh001_027_009+    i_027    tia_h_in_001_009+    14954.397020306033
Rh001_027_009-    i_027    tia_h_in_001_009-    14572.913754664809
Rh001_028_009+    i_028    tia_h_in_001_009+    14358.240407025502
Rh001_028_009-    i_028    tia_h_in_001_009-    14895.920038958528
Rh001_029_009+    i_029    tia_h_in_001_009+    14495.655236240435
Rh001_029_009-    i_029    tia_h_in_001_009-    14912.750356549494
Rh001_030_009+    i_030    tia_h_in_001_009+    14294.90103365636
Rh001_030_009-    i_030    tia_h_in_001_009-    15085.334031825856
Rh001_031_009+    i_031    tia_h_in_001_009+    13758.593693439454
Rh001_031_009-    i_031    tia_h_in_001_009-    14902.17938848914
Rh001_032_009+    i_032    tia_h_in_001_009+    12907.616358471982
Rh001_032_009-    i_032    tia_h_in_001_009-    14993.791518494725
Rh001_033_009+    i_033    tia_h_in_001_009+    12567.178920452216
Rh001_033_009-    i_033    tia_h_in_001_009-    14972.936847316132
Rh001_034_009+    i_034    tia_h_in_001_009+    14022.06329633376
Rh001_034_009-    i_034    tia_h_in_001_009-    14973.93503458376
Rh001_035_009+    i_035    tia_h_in_001_009+    14943.425198741255
Rh001_035_009-    i_035    tia_h_in_001_009-    13832.231701723675
Rh001_036_009+    i_036    tia_h_in_001_009+    14658.836006999456
Rh001_036_009-    i_036    tia_h_in_001_009-    14994.089003100422
Rh001_037_009+    i_037    tia_h_in_001_009+    14796.655884444348
Rh001_037_009-    i_037    tia_h_in_001_009-    14753.514825213113
Rh001_038_009+    i_038    tia_h_in_001_009+    15000
Rh001_038_009-    i_038    tia_h_in_001_009-    14972.651257198566
Rh001_039_009+    i_039    tia_h_in_001_009+    15099.243106519301
Rh001_039_009-    i_039    tia_h_in_001_009-    5000
Rh001_040_009+    i_040    tia_h_in_001_009+    13350.60150256076
Rh001_040_009-    i_040    tia_h_in_001_009-    14938.955580982296
Rh001_041_009+    i_041    tia_h_in_001_009+    12327.913481429552
Rh001_041_009-    i_041    tia_h_in_001_009-    14932.866278505431
Rh001_042_009+    i_042    tia_h_in_001_009+    14512.914965512457
Rh001_042_009-    i_042    tia_h_in_001_009-    14868.79065493288
Rh001_043_009+    i_043    tia_h_in_001_009+    14343.864025085468
Rh001_043_009-    i_043    tia_h_in_001_009-    15089.611146147881
Rh001_044_009+    i_044    tia_h_in_001_009+    12527.755733416383
Rh001_044_009-    i_044    tia_h_in_001_009-    14911.741111623962
Rh001_045_009+    i_045    tia_h_in_001_009+    12283.062676949197
Rh001_045_009-    i_045    tia_h_in_001_009-    15218.451008148239
Rh001_046_009+    i_046    tia_h_in_001_009+    14298.732495099779
Rh001_046_009-    i_046    tia_h_in_001_009-    14912.260794826429
Rh001_047_009+    i_047    tia_h_in_001_009+    12742.43178893808
Rh001_047_009-    i_047    tia_h_in_001_009-    5000
Rh001_048_009+    i_048    tia_h_in_001_009+    11101.4982674638
Rh001_048_009-    i_048    tia_h_in_001_009-    14954.306987911188
Rh001_049_009+    i_049    tia_h_in_001_009+    15091.877459083953
Rh001_049_009-    i_049    tia_h_in_001_009-    14602.656948678708
Rh001_050_009+    i_050    tia_h_in_001_009+    14371.068110715263
Rh001_050_009-    i_050    tia_h_in_001_009-    15086.04108869843
Rh001_051_009+    i_051    tia_h_in_001_009+    15036.967939666978
Rh001_051_009-    i_051    tia_h_in_001_009-    12586.058447200698
Rh001_052_009+    i_052    tia_h_in_001_009+    15000
Rh001_052_009-    i_052    tia_h_in_001_009-    14384.650985214568
Rh001_053_009+    i_053    tia_h_in_001_009+    5000
Rh001_053_009-    i_053    tia_h_in_001_009-    13502.495797275911
Rh001_054_009+    i_054    tia_h_in_001_009+    15132.935524399794
Rh001_054_009-    i_054    tia_h_in_001_009-    15119.86672750907
Rh001_055_009+    i_055    tia_h_in_001_009+    13360.042441061663
Rh001_055_009-    i_055    tia_h_in_001_009-    14994.349491232764
Rh001_056_009+    i_056    tia_h_in_001_009+    14911.33382003542
Rh001_056_009-    i_056    tia_h_in_001_009-    13081.089798102434
Rh001_057_009+    i_057    tia_h_in_001_009+    14942.253772367607
Rh001_057_009-    i_057    tia_h_in_001_009-    13574.25078274079
Rh001_058_009+    i_058    tia_h_in_001_009+    14903.560405937544
Rh001_058_009-    i_058    tia_h_in_001_009-    13342.147549746454
Rh001_059_009+    i_059    tia_h_in_001_009+    14349.71913263724
Rh001_059_009-    i_059    tia_h_in_001_009-    14930.749471777757
Rh001_060_009+    i_060    tia_h_in_001_009+    14982.180447162222
Rh001_060_009-    i_060    tia_h_in_001_009-    13188.372240241528
Rh001_061_009+    i_061    tia_h_in_001_009+    15223.153700226405
Rh001_061_009-    i_061    tia_h_in_001_009-    12651.181347181566
Rh001_062_009+    i_062    tia_h_in_001_009+    14955.43964940503
Rh001_062_009-    i_062    tia_h_in_001_009-    13554.98282464362
Rh001_063_009+    i_063    tia_h_in_001_009+    15048.70919560666
Rh001_063_009-    i_063    tia_h_in_001_009-    10514.43757108437
Rh001_064_009+    i_064    tia_h_in_001_009+    14921.451246296649
Rh001_064_009-    i_064    tia_h_in_001_009-    9234.391180576773

* Neuron 10
Rh001_001_010+    i_001    tia_h_in_001_010+    14104.440096040522
Rh001_001_010-    i_001    tia_h_in_001_010-    14959.656964314137
Rh001_002_010+    i_002    tia_h_in_001_010+    14962.70031579976
Rh001_002_010-    i_002    tia_h_in_001_010-    13787.390183937405
Rh001_003_010+    i_003    tia_h_in_001_010+    14788.000232186827
Rh001_003_010-    i_003    tia_h_in_001_010-    15157.882239431505
Rh001_004_010+    i_004    tia_h_in_001_010+    13677.260154285967
Rh001_004_010-    i_004    tia_h_in_001_010-    14747.786964677462
Rh001_005_010+    i_005    tia_h_in_001_010+    14738.319831853587
Rh001_005_010-    i_005    tia_h_in_001_010-    14838.918495720101
Rh001_006_010+    i_006    tia_h_in_001_010+    14666.852467904002
Rh001_006_010-    i_006    tia_h_in_001_010-    15079.760700371571
Rh001_007_010+    i_007    tia_h_in_001_010+    14832.398332260382
Rh001_007_010-    i_007    tia_h_in_001_010-    13964.678635298447
Rh001_008_010+    i_008    tia_h_in_001_010+    14975.845922169901
Rh001_008_010-    i_008    tia_h_in_001_010-    14906.555689985262
Rh001_009_010+    i_009    tia_h_in_001_010+    15173.72285575836
Rh001_009_010-    i_009    tia_h_in_001_010-    14954.69446293566
Rh001_010_010+    i_010    tia_h_in_001_010+    14520.344001545958
Rh001_010_010-    i_010    tia_h_in_001_010-    15055.020518977346
Rh001_011_010+    i_011    tia_h_in_001_010+    5000
Rh001_011_010-    i_011    tia_h_in_001_010-    15149.795277668447
Rh001_012_010+    i_012    tia_h_in_001_010+    13829.367810336396
Rh001_012_010-    i_012    tia_h_in_001_010-    14927.147978440325
Rh001_013_010+    i_013    tia_h_in_001_010+    15036.2538469854
Rh001_013_010-    i_013    tia_h_in_001_010-    13846.99926202397
Rh001_014_010+    i_014    tia_h_in_001_010+    5000
Rh001_014_010-    i_014    tia_h_in_001_010-    15075.176822782512
Rh001_015_010+    i_015    tia_h_in_001_010+    14772.279482943257
Rh001_015_010-    i_015    tia_h_in_001_010-    15000
Rh001_016_010+    i_016    tia_h_in_001_010+    15093.347214591866
Rh001_016_010-    i_016    tia_h_in_001_010-    13808.69655510535
Rh001_017_010+    i_017    tia_h_in_001_010+    15104.980947182761
Rh001_017_010-    i_017    tia_h_in_001_010-    14773.389900691283
Rh001_018_010+    i_018    tia_h_in_001_010+    14999.82924464292
Rh001_018_010-    i_018    tia_h_in_001_010-    13666.04034534899
Rh001_019_010+    i_019    tia_h_in_001_010+    14291.008662318542
Rh001_019_010-    i_019    tia_h_in_001_010-    15037.352937475498
Rh001_020_010+    i_020    tia_h_in_001_010+    14884.482947243177
Rh001_020_010-    i_020    tia_h_in_001_010-    14974.999489362015
Rh001_021_010+    i_021    tia_h_in_001_010+    14864.94185898948
Rh001_021_010-    i_021    tia_h_in_001_010-    14091.609874239379
Rh001_022_010+    i_022    tia_h_in_001_010+    14101.71647924013
Rh001_022_010-    i_022    tia_h_in_001_010-    15071.507614096754
Rh001_023_010+    i_023    tia_h_in_001_010+    5000
Rh001_023_010-    i_023    tia_h_in_001_010-    13475.017257336127
Rh001_024_010+    i_024    tia_h_in_001_010+    14907.16147222661
Rh001_024_010-    i_024    tia_h_in_001_010-    14274.262524904365
Rh001_025_010+    i_025    tia_h_in_001_010+    15186.993763571207
Rh001_025_010-    i_025    tia_h_in_001_010-    14475.75439024654
Rh001_026_010+    i_026    tia_h_in_001_010+    15130.129615564478
Rh001_026_010-    i_026    tia_h_in_001_010-    13718.605209606774
Rh001_027_010+    i_027    tia_h_in_001_010+    5000
Rh001_027_010-    i_027    tia_h_in_001_010-    13755.004717489826
Rh001_028_010+    i_028    tia_h_in_001_010+    5000
Rh001_028_010-    i_028    tia_h_in_001_010-    14840.019476560996
Rh001_029_010+    i_029    tia_h_in_001_010+    5000
Rh001_029_010-    i_029    tia_h_in_001_010-    15011.155597151082
Rh001_030_010+    i_030    tia_h_in_001_010+    13701.307819144566
Rh001_030_010-    i_030    tia_h_in_001_010-    15010.278493547301
Rh001_031_010+    i_031    tia_h_in_001_010+    15000
Rh001_031_010-    i_031    tia_h_in_001_010-    15034.204246281564
Rh001_032_010+    i_032    tia_h_in_001_010+    14872.529066164398
Rh001_032_010-    i_032    tia_h_in_001_010-    14026.720545228198
Rh001_033_010+    i_033    tia_h_in_001_010+    15196.10976442988
Rh001_033_010-    i_033    tia_h_in_001_010-    13836.75319404518
Rh001_034_010+    i_034    tia_h_in_001_010+    13722.10398718929
Rh001_034_010-    i_034    tia_h_in_001_010-    14870.765608214966
Rh001_035_010+    i_035    tia_h_in_001_010+    14550.666347684726
Rh001_035_010-    i_035    tia_h_in_001_010-    15112.715344659186
Rh001_036_010+    i_036    tia_h_in_001_010+    14980.474567549487
Rh001_036_010-    i_036    tia_h_in_001_010-    14978.424072740803
Rh001_037_010+    i_037    tia_h_in_001_010+    14626.412225495518
Rh001_037_010-    i_037    tia_h_in_001_010-    15267.28964996313
Rh001_038_010+    i_038    tia_h_in_001_010+    14979.968559677154
Rh001_038_010-    i_038    tia_h_in_001_010-    13879.358398918825
Rh001_039_010+    i_039    tia_h_in_001_010+    15162.311786790344
Rh001_039_010-    i_039    tia_h_in_001_010-    5000
Rh001_040_010+    i_040    tia_h_in_001_010+    13791.633791788936
Rh001_040_010-    i_040    tia_h_in_001_010-    15080.4524272124
Rh001_041_010+    i_041    tia_h_in_001_010+    15000
Rh001_041_010-    i_041    tia_h_in_001_010-    14625.056480247425
Rh001_042_010+    i_042    tia_h_in_001_010+    14925.236943222386
Rh001_042_010-    i_042    tia_h_in_001_010-    14884.736907852157
Rh001_043_010+    i_043    tia_h_in_001_010+    14938.527740555593
Rh001_043_010-    i_043    tia_h_in_001_010-    13850.597127872494
Rh001_044_010+    i_044    tia_h_in_001_010+    15226.56994458086
Rh001_044_010-    i_044    tia_h_in_001_010-    14113.708858494372
Rh001_045_010+    i_045    tia_h_in_001_010+    15078.708776604552
Rh001_045_010-    i_045    tia_h_in_001_010-    14888.692698323977
Rh001_046_010+    i_046    tia_h_in_001_010+    15141.854382862402
Rh001_046_010-    i_046    tia_h_in_001_010-    13922.965942778323
Rh001_047_010+    i_047    tia_h_in_001_010+    15207.56982372236
Rh001_047_010-    i_047    tia_h_in_001_010-    14926.921820937543
Rh001_048_010+    i_048    tia_h_in_001_010+    14446.404543789411
Rh001_048_010-    i_048    tia_h_in_001_010-    15041.869460637516
Rh001_049_010+    i_049    tia_h_in_001_010+    5000
Rh001_049_010-    i_049    tia_h_in_001_010-    13504.338689543196
Rh001_050_010+    i_050    tia_h_in_001_010+    14669.221775591923
Rh001_050_010-    i_050    tia_h_in_001_010-    15038.728330997705
Rh001_051_010+    i_051    tia_h_in_001_010+    14838.95176536625
Rh001_051_010-    i_051    tia_h_in_001_010-    13961.117129585413
Rh001_052_010+    i_052    tia_h_in_001_010+    15145.040315725384
Rh001_052_010-    i_052    tia_h_in_001_010-    14239.915112615148
Rh001_053_010+    i_053    tia_h_in_001_010+    15000
Rh001_053_010-    i_053    tia_h_in_001_010-    14863.128110478408
Rh001_054_010+    i_054    tia_h_in_001_010+    13852.635858660213
Rh001_054_010-    i_054    tia_h_in_001_010-    5000
Rh001_055_010+    i_055    tia_h_in_001_010+    15110.772608799438
Rh001_055_010-    i_055    tia_h_in_001_010-    14233.515713120216
Rh001_056_010+    i_056    tia_h_in_001_010+    14870.76164937791
Rh001_056_010-    i_056    tia_h_in_001_010-    14318.497817398696
Rh001_057_010+    i_057    tia_h_in_001_010+    14949.600606587079
Rh001_057_010-    i_057    tia_h_in_001_010-    13728.86367341189
Rh001_058_010+    i_058    tia_h_in_001_010+    5000
Rh001_058_010-    i_058    tia_h_in_001_010-    5000
Rh001_059_010+    i_059    tia_h_in_001_010+    14929.735195658
Rh001_059_010-    i_059    tia_h_in_001_010-    13731.01600714326
Rh001_060_010+    i_060    tia_h_in_001_010+    15151.328520633013
Rh001_060_010-    i_060    tia_h_in_001_010-    14484.7908590058
Rh001_061_010+    i_061    tia_h_in_001_010+    14849.812905365285
Rh001_061_010-    i_061    tia_h_in_001_010-    14988.889685724816
Rh001_062_010+    i_062    tia_h_in_001_010+    15245.026785884616
Rh001_062_010-    i_062    tia_h_in_001_010-    13569.845775389822
Rh001_063_010+    i_063    tia_h_in_001_010+    13658.036527951499
Rh001_063_010-    i_063    tia_h_in_001_010-    15040.622173539632
Rh001_064_010+    i_064    tia_h_in_001_010+    14210.298783855278
Rh001_064_010-    i_064    tia_h_in_001_010-    15337.638024215456

* Neuron 11
Rh001_001_011+    i_001    tia_h_in_001_011+    14944.068053355328
Rh001_001_011-    i_001    tia_h_in_001_011-    9397.832733013933
Rh001_002_011+    i_002    tia_h_in_001_011+    15145.586467300922
Rh001_002_011-    i_002    tia_h_in_001_011-    11654.361842859797
Rh001_003_011+    i_003    tia_h_in_001_011+    15156.876650350232
Rh001_003_011-    i_003    tia_h_in_001_011-    11930.574362814223
Rh001_004_011+    i_004    tia_h_in_001_011+    14795.895073604597
Rh001_004_011-    i_004    tia_h_in_001_011-    11503.720200673357
Rh001_005_011+    i_005    tia_h_in_001_011+    14797.117476018706
Rh001_005_011-    i_005    tia_h_in_001_011-    12405.974392980437
Rh001_006_011+    i_006    tia_h_in_001_011+    15010.294527655415
Rh001_006_011-    i_006    tia_h_in_001_011-    11796.07759215735
Rh001_007_011+    i_007    tia_h_in_001_011+    14388.44464080808
Rh001_007_011-    i_007    tia_h_in_001_011-    5000
Rh001_008_011+    i_008    tia_h_in_001_011+    14905.985173996625
Rh001_008_011-    i_008    tia_h_in_001_011-    14624.245905752085
Rh001_009_011+    i_009    tia_h_in_001_011+    12723.37444619866
Rh001_009_011-    i_009    tia_h_in_001_011-    14867.945458713672
Rh001_010_011+    i_010    tia_h_in_001_011+    12842.030373731463
Rh001_010_011-    i_010    tia_h_in_001_011-    14945.50019123117
Rh001_011_011+    i_011    tia_h_in_001_011+    15000
Rh001_011_011-    i_011    tia_h_in_001_011-    15042.91744323779
Rh001_012_011+    i_012    tia_h_in_001_011+    12303.152897054471
Rh001_012_011-    i_012    tia_h_in_001_011-    15027.558505185225
Rh001_013_011+    i_013    tia_h_in_001_011+    14112.11725859992
Rh001_013_011-    i_013    tia_h_in_001_011-    14742.085109833095
Rh001_014_011+    i_014    tia_h_in_001_011+    15325.006603296159
Rh001_014_011-    i_014    tia_h_in_001_011-    14479.461362210819
Rh001_015_011+    i_015    tia_h_in_001_011+    15055.727968530899
Rh001_015_011-    i_015    tia_h_in_001_011-    13759.666333974901
Rh001_016_011+    i_016    tia_h_in_001_011+    15000
Rh001_016_011-    i_016    tia_h_in_001_011-    14103.95720581825
Rh001_017_011+    i_017    tia_h_in_001_011+    12659.654050975552
Rh001_017_011-    i_017    tia_h_in_001_011-    14888.85608391504
Rh001_018_011+    i_018    tia_h_in_001_011+    12574.251219716223
Rh001_018_011-    i_018    tia_h_in_001_011-    15184.440457760982
Rh001_019_011+    i_019    tia_h_in_001_011+    15144.966712752068
Rh001_019_011-    i_019    tia_h_in_001_011-    13684.405770760375
Rh001_020_011+    i_020    tia_h_in_001_011+    12971.540788900742
Rh001_020_011-    i_020    tia_h_in_001_011-    14793.930156487539
Rh001_021_011+    i_021    tia_h_in_001_011+    11592.290338253613
Rh001_021_011-    i_021    tia_h_in_001_011-    15086.742157930337
Rh001_022_011+    i_022    tia_h_in_001_011+    14054.892298082415
Rh001_022_011-    i_022    tia_h_in_001_011-    15116.23374685622
Rh001_023_011+    i_023    tia_h_in_001_011+    14926.511830034346
Rh001_023_011-    i_023    tia_h_in_001_011-    14805.344779664514
Rh001_024_011+    i_024    tia_h_in_001_011+    14538.565079922057
Rh001_024_011-    i_024    tia_h_in_001_011-    14695.66204334603
Rh001_025_011+    i_025    tia_h_in_001_011+    13448.71433168322
Rh001_025_011-    i_025    tia_h_in_001_011-    15000
Rh001_026_011+    i_026    tia_h_in_001_011+    15018.198368873407
Rh001_026_011-    i_026    tia_h_in_001_011-    15000
Rh001_027_011+    i_027    tia_h_in_001_011+    15000
Rh001_027_011-    i_027    tia_h_in_001_011-    14840.98064808545
Rh001_028_011+    i_028    tia_h_in_001_011+    14159.63206409672
Rh001_028_011-    i_028    tia_h_in_001_011-    15050.796661034943
Rh001_029_011+    i_029    tia_h_in_001_011+    14502.726278610213
Rh001_029_011-    i_029    tia_h_in_001_011-    15043.692481548107
Rh001_030_011+    i_030    tia_h_in_001_011+    14213.264776050373
Rh001_030_011-    i_030    tia_h_in_001_011-    15111.117977130934
Rh001_031_011+    i_031    tia_h_in_001_011+    13439.46483649989
Rh001_031_011-    i_031    tia_h_in_001_011-    15004.241401349158
Rh001_032_011+    i_032    tia_h_in_001_011+    14161.289290532863
Rh001_032_011-    i_032    tia_h_in_001_011-    5000
Rh001_033_011+    i_033    tia_h_in_001_011+    15007.301470503127
Rh001_033_011-    i_033    tia_h_in_001_011-    14828.839223118412
Rh001_034_011+    i_034    tia_h_in_001_011+    15000
Rh001_034_011-    i_034    tia_h_in_001_011-    14927.22288248517
Rh001_035_011+    i_035    tia_h_in_001_011+    5000
Rh001_035_011-    i_035    tia_h_in_001_011-    14916.383770196604
Rh001_036_011+    i_036    tia_h_in_001_011+    14970.87931365518
Rh001_036_011-    i_036    tia_h_in_001_011-    12224.533135323496
Rh001_037_011+    i_037    tia_h_in_001_011+    15138.162637851712
Rh001_037_011-    i_037    tia_h_in_001_011-    14928.242078221292
Rh001_038_011+    i_038    tia_h_in_001_011+    13802.875247830683
Rh001_038_011-    i_038    tia_h_in_001_011-    5000
Rh001_039_011+    i_039    tia_h_in_001_011+    13718.715564642232
Rh001_039_011-    i_039    tia_h_in_001_011-    14979.98164161206
Rh001_040_011+    i_040    tia_h_in_001_011+    15000
Rh001_040_011-    i_040    tia_h_in_001_011-    12714.779320903202
Rh001_041_011+    i_041    tia_h_in_001_011+    14286.123504328467
Rh001_041_011-    i_041    tia_h_in_001_011-    14914.502139963715
Rh001_042_011+    i_042    tia_h_in_001_011+    15064.267104882632
Rh001_042_011-    i_042    tia_h_in_001_011-    14812.390675281335
Rh001_043_011+    i_043    tia_h_in_001_011+    15115.88295906487
Rh001_043_011-    i_043    tia_h_in_001_011-    12987.725892945837
Rh001_044_011+    i_044    tia_h_in_001_011+    14923.890710901862
Rh001_044_011-    i_044    tia_h_in_001_011-    13306.988103026266
Rh001_045_011+    i_045    tia_h_in_001_011+    14890.062424602767
Rh001_045_011-    i_045    tia_h_in_001_011-    12202.4792643043
Rh001_046_011+    i_046    tia_h_in_001_011+    15008.015623423293
Rh001_046_011-    i_046    tia_h_in_001_011-    13459.077542034207
Rh001_047_011+    i_047    tia_h_in_001_011+    13673.59483762776
Rh001_047_011-    i_047    tia_h_in_001_011-    14972.978136737534
Rh001_048_011+    i_048    tia_h_in_001_011+    14949.57347222813
Rh001_048_011-    i_048    tia_h_in_001_011-    5000
Rh001_049_011+    i_049    tia_h_in_001_011+    14962.361306836865
Rh001_049_011-    i_049    tia_h_in_001_011-    13925.41568622554
Rh001_050_011+    i_050    tia_h_in_001_011+    14059.403330679397
Rh001_050_011-    i_050    tia_h_in_001_011-    15068.693289292733
Rh001_051_011+    i_051    tia_h_in_001_011+    14134.24936047129
Rh001_051_011-    i_051    tia_h_in_001_011-    15052.380389954094
Rh001_052_011+    i_052    tia_h_in_001_011+    15000
Rh001_052_011-    i_052    tia_h_in_001_011-    15205.83597495004
Rh001_053_011+    i_053    tia_h_in_001_011+    13327.937974433766
Rh001_053_011-    i_053    tia_h_in_001_011-    14733.846655722175
Rh001_054_011+    i_054    tia_h_in_001_011+    5000
Rh001_054_011-    i_054    tia_h_in_001_011-    14249.309667461257
Rh001_055_011+    i_055    tia_h_in_001_011+    14905.391011077183
Rh001_055_011-    i_055    tia_h_in_001_011-    12300.895289499766
Rh001_056_011+    i_056    tia_h_in_001_011+    13826.105638566156
Rh001_056_011-    i_056    tia_h_in_001_011-    14946.5716694169
Rh001_057_011+    i_057    tia_h_in_001_011+    14332.205237429984
Rh001_057_011-    i_057    tia_h_in_001_011-    14832.579105480907
Rh001_058_011+    i_058    tia_h_in_001_011+    14933.905416381609
Rh001_058_011-    i_058    tia_h_in_001_011-    14702.472210298027
Rh001_059_011+    i_059    tia_h_in_001_011+    13375.740304774341
Rh001_059_011-    i_059    tia_h_in_001_011-    14854.796860661827
Rh001_060_011+    i_060    tia_h_in_001_011+    15003.019579112732
Rh001_060_011-    i_060    tia_h_in_001_011-    14786.89953031748
Rh001_061_011+    i_061    tia_h_in_001_011+    14072.115824530616
Rh001_061_011-    i_061    tia_h_in_001_011-    14938.130157524305
Rh001_062_011+    i_062    tia_h_in_001_011+    14825.5983706507
Rh001_062_011-    i_062    tia_h_in_001_011-    14507.450300567963
Rh001_063_011+    i_063    tia_h_in_001_011+    12641.992244907573
Rh001_063_011-    i_063    tia_h_in_001_011-    15093.780899258847
Rh001_064_011+    i_064    tia_h_in_001_011+    15077.756419880867
Rh001_064_011-    i_064    tia_h_in_001_011-    14830.874356117021

* Neuron 12
Rh001_001_012+    i_001    tia_h_in_001_012+    15048.794992820045
Rh001_001_012-    i_001    tia_h_in_001_012-    11872.280684646543
Rh001_002_012+    i_002    tia_h_in_001_012+    15000
Rh001_002_012-    i_002    tia_h_in_001_012-    15000
Rh001_003_012+    i_003    tia_h_in_001_012+    5000
Rh001_003_012-    i_003    tia_h_in_001_012-    11970.598978000498
Rh001_004_012+    i_004    tia_h_in_001_012+    15000
Rh001_004_012-    i_004    tia_h_in_001_012-    5000
Rh001_005_012+    i_005    tia_h_in_001_012+    13711.18010727793
Rh001_005_012-    i_005    tia_h_in_001_012-    15084.45397756932
Rh001_006_012+    i_006    tia_h_in_001_012+    15000
Rh001_006_012-    i_006    tia_h_in_001_012-    13361.086982633904
Rh001_007_012+    i_007    tia_h_in_001_012+    14983.04007833722
Rh001_007_012-    i_007    tia_h_in_001_012-    14969.510709765224
Rh001_008_012+    i_008    tia_h_in_001_012+    15000
Rh001_008_012-    i_008    tia_h_in_001_012-    14708.371296546848
Rh001_009_012+    i_009    tia_h_in_001_012+    14658.040021397928
Rh001_009_012-    i_009    tia_h_in_001_012-    5000
Rh001_010_012+    i_010    tia_h_in_001_012+    5000
Rh001_010_012-    i_010    tia_h_in_001_012-    12165.129785721036
Rh001_011_012+    i_011    tia_h_in_001_012+    15033.324644391252
Rh001_011_012-    i_011    tia_h_in_001_012-    13629.967618294731
Rh001_012_012+    i_012    tia_h_in_001_012+    15223.621775691834
Rh001_012_012-    i_012    tia_h_in_001_012-    12417.384140152282
Rh001_013_012+    i_013    tia_h_in_001_012+    5000
Rh001_013_012-    i_013    tia_h_in_001_012-    14992.74728315838
Rh001_014_012+    i_014    tia_h_in_001_012+    13058.126798261852
Rh001_014_012-    i_014    tia_h_in_001_012-    14891.50558313948
Rh001_015_012+    i_015    tia_h_in_001_012+    14118.012109547959
Rh001_015_012-    i_015    tia_h_in_001_012-    14894.850692232218
Rh001_016_012+    i_016    tia_h_in_001_012+    14691.411306427926
Rh001_016_012-    i_016    tia_h_in_001_012-    14856.798950681456
Rh001_017_012+    i_017    tia_h_in_001_012+    15083.950960673486
Rh001_017_012-    i_017    tia_h_in_001_012-    13721.169198054196
Rh001_018_012+    i_018    tia_h_in_001_012+    12619.210326627695
Rh001_018_012-    i_018    tia_h_in_001_012-    15000
Rh001_019_012+    i_019    tia_h_in_001_012+    14370.133037281674
Rh001_019_012-    i_019    tia_h_in_001_012-    14905.550520308621
Rh001_020_012+    i_020    tia_h_in_001_012+    14968.353347475333
Rh001_020_012-    i_020    tia_h_in_001_012-    11415.173472066652
Rh001_021_012+    i_021    tia_h_in_001_012+    14948.378838430302
Rh001_021_012-    i_021    tia_h_in_001_012-    14341.67205460187
Rh001_022_012+    i_022    tia_h_in_001_012+    15126.419904929378
Rh001_022_012-    i_022    tia_h_in_001_012-    13472.715160065605
Rh001_023_012+    i_023    tia_h_in_001_012+    12750.665196454285
Rh001_023_012-    i_023    tia_h_in_001_012-    15078.519915506542
Rh001_024_012+    i_024    tia_h_in_001_012+    14927.827515641353
Rh001_024_012-    i_024    tia_h_in_001_012-    14440.992072550816
Rh001_025_012+    i_025    tia_h_in_001_012+    15050.658552257042
Rh001_025_012-    i_025    tia_h_in_001_012-    12737.146514377873
Rh001_026_012+    i_026    tia_h_in_001_012+    14335.26115147575
Rh001_026_012-    i_026    tia_h_in_001_012-    15242.148723735441
Rh001_027_012+    i_027    tia_h_in_001_012+    12683.508671264046
Rh001_027_012-    i_027    tia_h_in_001_012-    15172.842580868612
Rh001_028_012+    i_028    tia_h_in_001_012+    13640.963681686679
Rh001_028_012-    i_028    tia_h_in_001_012-    14947.772319178512
Rh001_029_012+    i_029    tia_h_in_001_012+    15149.27175959023
Rh001_029_012-    i_029    tia_h_in_001_012-    14279.402008469771
Rh001_030_012+    i_030    tia_h_in_001_012+    15000
Rh001_030_012-    i_030    tia_h_in_001_012-    14225.38910407424
Rh001_031_012+    i_031    tia_h_in_001_012+    13019.442826355025
Rh001_031_012-    i_031    tia_h_in_001_012-    15155.05510952078
Rh001_032_012+    i_032    tia_h_in_001_012+    11444.230804586565
Rh001_032_012-    i_032    tia_h_in_001_012-    14976.477351856216
Rh001_033_012+    i_033    tia_h_in_001_012+    12888.070503852674
Rh001_033_012-    i_033    tia_h_in_001_012-    15008.393593291017
Rh001_034_012+    i_034    tia_h_in_001_012+    15088.025562013923
Rh001_034_012-    i_034    tia_h_in_001_012-    15042.837472022347
Rh001_035_012+    i_035    tia_h_in_001_012+    13699.464928861045
Rh001_035_012-    i_035    tia_h_in_001_012-    15016.038244398755
Rh001_036_012+    i_036    tia_h_in_001_012+    15000
Rh001_036_012-    i_036    tia_h_in_001_012-    15049.762028909558
Rh001_037_012+    i_037    tia_h_in_001_012+    15000
Rh001_037_012-    i_037    tia_h_in_001_012-    14914.06476786967
Rh001_038_012+    i_038    tia_h_in_001_012+    14457.433691733335
Rh001_038_012-    i_038    tia_h_in_001_012-    15058.61736631762
Rh001_039_012+    i_039    tia_h_in_001_012+    13823.97591146832
Rh001_039_012-    i_039    tia_h_in_001_012-    15208.965222996407
Rh001_040_012+    i_040    tia_h_in_001_012+    14970.845706366646
Rh001_040_012-    i_040    tia_h_in_001_012-    13484.869671302531
Rh001_041_012+    i_041    tia_h_in_001_012+    12527.382345607837
Rh001_041_012-    i_041    tia_h_in_001_012-    15125.358026309648
Rh001_042_012+    i_042    tia_h_in_001_012+    13640.36815114336
Rh001_042_012-    i_042    tia_h_in_001_012-    14905.04687544724
Rh001_043_012+    i_043    tia_h_in_001_012+    14987.219450587017
Rh001_043_012-    i_043    tia_h_in_001_012-    15059.67685441664
Rh001_044_012+    i_044    tia_h_in_001_012+    15000
Rh001_044_012-    i_044    tia_h_in_001_012-    15187.228056759472
Rh001_045_012+    i_045    tia_h_in_001_012+    14922.299830879609
Rh001_045_012-    i_045    tia_h_in_001_012-    13237.422432000028
Rh001_046_012+    i_046    tia_h_in_001_012+    5000
Rh001_046_012-    i_046    tia_h_in_001_012-    12910.457250715495
Rh001_047_012+    i_047    tia_h_in_001_012+    14258.57332555383
Rh001_047_012-    i_047    tia_h_in_001_012-    14916.961896466217
Rh001_048_012+    i_048    tia_h_in_001_012+    15122.311818879363
Rh001_048_012-    i_048    tia_h_in_001_012-    12825.129871151483
Rh001_049_012+    i_049    tia_h_in_001_012+    12943.219053572453
Rh001_049_012-    i_049    tia_h_in_001_012-    15156.528409944129
Rh001_050_012+    i_050    tia_h_in_001_012+    15000
Rh001_050_012-    i_050    tia_h_in_001_012-    15000
Rh001_051_012+    i_051    tia_h_in_001_012+    15014.357307757442
Rh001_051_012-    i_051    tia_h_in_001_012-    14410.43561110768
Rh001_052_012+    i_052    tia_h_in_001_012+    14403.556100362619
Rh001_052_012-    i_052    tia_h_in_001_012-    15018.608134979584
Rh001_053_012+    i_053    tia_h_in_001_012+    5000
Rh001_053_012-    i_053    tia_h_in_001_012-    14918.052325604738
Rh001_054_012+    i_054    tia_h_in_001_012+    14097.902582092725
Rh001_054_012-    i_054    tia_h_in_001_012-    15192.468372818694
Rh001_055_012+    i_055    tia_h_in_001_012+    15000
Rh001_055_012-    i_055    tia_h_in_001_012-    13067.572475290555
Rh001_056_012+    i_056    tia_h_in_001_012+    14949.686984389611
Rh001_056_012-    i_056    tia_h_in_001_012-    15044.700658043997
Rh001_057_012+    i_057    tia_h_in_001_012+    14888.928119919763
Rh001_057_012-    i_057    tia_h_in_001_012-    12987.356108265305
Rh001_058_012+    i_058    tia_h_in_001_012+    14696.234861686822
Rh001_058_012-    i_058    tia_h_in_001_012-    15096.004230731869
Rh001_059_012+    i_059    tia_h_in_001_012+    15008.550734060476
Rh001_059_012-    i_059    tia_h_in_001_012-    13316.843320984563
Rh001_060_012+    i_060    tia_h_in_001_012+    15042.390887666073
Rh001_060_012-    i_060    tia_h_in_001_012-    13186.467796626346
Rh001_061_012+    i_061    tia_h_in_001_012+    13988.287540636498
Rh001_061_012-    i_061    tia_h_in_001_012-    15133.6630035466
Rh001_062_012+    i_062    tia_h_in_001_012+    15000
Rh001_062_012-    i_062    tia_h_in_001_012-    12837.426806966261
Rh001_063_012+    i_063    tia_h_in_001_012+    15090.500656219343
Rh001_063_012-    i_063    tia_h_in_001_012-    15000
Rh001_064_012+    i_064    tia_h_in_001_012+    15186.886280045457
Rh001_064_012-    i_064    tia_h_in_001_012-    13672.561792002025

* Neuron 13
Rh001_001_013+    i_001    tia_h_in_001_013+    15086.553149342275
Rh001_001_013-    i_001    tia_h_in_001_013-    5000
Rh001_002_013+    i_002    tia_h_in_001_013+    15197.571927601575
Rh001_002_013-    i_002    tia_h_in_001_013-    9793.000599289424
Rh001_003_013+    i_003    tia_h_in_001_013+    15102.488885007351
Rh001_003_013-    i_003    tia_h_in_001_013-    12277.550464621601
Rh001_004_013+    i_004    tia_h_in_001_013+    15128.780351956815
Rh001_004_013-    i_004    tia_h_in_001_013-    12490.797595998078
Rh001_005_013+    i_005    tia_h_in_001_013+    15154.9973916995
Rh001_005_013-    i_005    tia_h_in_001_013-    5000
Rh001_006_013+    i_006    tia_h_in_001_013+    13306.802324145427
Rh001_006_013-    i_006    tia_h_in_001_013-    5000
Rh001_007_013+    i_007    tia_h_in_001_013+    5000
Rh001_007_013-    i_007    tia_h_in_001_013-    13655.530289638156
Rh001_008_013+    i_008    tia_h_in_001_013+    13831.037095458174
Rh001_008_013-    i_008    tia_h_in_001_013-    15087.674839405994
Rh001_009_013+    i_009    tia_h_in_001_013+    14214.716345722574
Rh001_009_013-    i_009    tia_h_in_001_013-    14848.466301058608
Rh001_010_013+    i_010    tia_h_in_001_013+    15000
Rh001_010_013-    i_010    tia_h_in_001_013-    15102.279044463887
Rh001_011_013+    i_011    tia_h_in_001_013+    13014.242779287164
Rh001_011_013-    i_011    tia_h_in_001_013-    14894.996070858522
Rh001_012_013+    i_012    tia_h_in_001_013+    15061.556279687595
Rh001_012_013-    i_012    tia_h_in_001_013-    13760.57790393979
Rh001_013_013+    i_013    tia_h_in_001_013+    5000
Rh001_013_013-    i_013    tia_h_in_001_013-    14976.617682186614
Rh001_014_013+    i_014    tia_h_in_001_013+    14959.954279365467
Rh001_014_013-    i_014    tia_h_in_001_013-    13552.438375543165
Rh001_015_013+    i_015    tia_h_in_001_013+    14741.33934493659
Rh001_015_013-    i_015    tia_h_in_001_013-    15095.339024337214
Rh001_016_013+    i_016    tia_h_in_001_013+    14218.133542370077
Rh001_016_013-    i_016    tia_h_in_001_013-    14863.327153801289
Rh001_017_013+    i_017    tia_h_in_001_013+    10794.035400135424
Rh001_017_013-    i_017    tia_h_in_001_013-    14962.595122868091
Rh001_018_013+    i_018    tia_h_in_001_013+    12593.03981604596
Rh001_018_013-    i_018    tia_h_in_001_013-    15044.710478094967
Rh001_019_013+    i_019    tia_h_in_001_013+    12854.143955439222
Rh001_019_013-    i_019    tia_h_in_001_013-    15176.861405104462
Rh001_020_013+    i_020    tia_h_in_001_013+    14624.971963743268
Rh001_020_013-    i_020    tia_h_in_001_013-    15046.821496694889
Rh001_021_013+    i_021    tia_h_in_001_013+    14728.572730078607
Rh001_021_013-    i_021    tia_h_in_001_013-    13963.547024318357
Rh001_022_013+    i_022    tia_h_in_001_013+    14812.227108607845
Rh001_022_013-    i_022    tia_h_in_001_013-    13866.883948440629
Rh001_023_013+    i_023    tia_h_in_001_013+    14944.15980615354
Rh001_023_013-    i_023    tia_h_in_001_013-    13107.286825035664
Rh001_024_013+    i_024    tia_h_in_001_013+    15040.268199808446
Rh001_024_013-    i_024    tia_h_in_001_013-    11819.99249599306
Rh001_025_013+    i_025    tia_h_in_001_013+    5000
Rh001_025_013-    i_025    tia_h_in_001_013-    14951.398569322228
Rh001_026_013+    i_026    tia_h_in_001_013+    13942.847169832537
Rh001_026_013-    i_026    tia_h_in_001_013-    15080.796213463573
Rh001_027_013+    i_027    tia_h_in_001_013+    13302.032452774132
Rh001_027_013-    i_027    tia_h_in_001_013-    14933.7197228962
Rh001_028_013+    i_028    tia_h_in_001_013+    15000
Rh001_028_013-    i_028    tia_h_in_001_013-    5000
Rh001_029_013+    i_029    tia_h_in_001_013+    14909.707384197116
Rh001_029_013-    i_029    tia_h_in_001_013-    12455.783716527902
Rh001_030_013+    i_030    tia_h_in_001_013+    13857.977267205297
Rh001_030_013-    i_030    tia_h_in_001_013-    5000
Rh001_031_013+    i_031    tia_h_in_001_013+    14929.339455569847
Rh001_031_013-    i_031    tia_h_in_001_013-    14125.60833335076
Rh001_032_013+    i_032    tia_h_in_001_013+    14123.0765480127
Rh001_032_013-    i_032    tia_h_in_001_013-    14987.349679577756
Rh001_033_013+    i_033    tia_h_in_001_013+    5000
Rh001_033_013-    i_033    tia_h_in_001_013-    14288.2254760844
Rh001_034_013+    i_034    tia_h_in_001_013+    15026.201738330248
Rh001_034_013-    i_034    tia_h_in_001_013-    13865.109932451069
Rh001_035_013+    i_035    tia_h_in_001_013+    15024.176460809556
Rh001_035_013-    i_035    tia_h_in_001_013-    14646.686990694554
Rh001_036_013+    i_036    tia_h_in_001_013+    5000
Rh001_036_013-    i_036    tia_h_in_001_013-    5000
Rh001_037_013+    i_037    tia_h_in_001_013+    12114.281822250017
Rh001_037_013-    i_037    tia_h_in_001_013-    14873.786731265076
Rh001_038_013+    i_038    tia_h_in_001_013+    5000
Rh001_038_013-    i_038    tia_h_in_001_013-    15000
Rh001_039_013+    i_039    tia_h_in_001_013+    15000
Rh001_039_013-    i_039    tia_h_in_001_013-    15113.73577731236
Rh001_040_013+    i_040    tia_h_in_001_013+    15128.979487209877
Rh001_040_013-    i_040    tia_h_in_001_013-    13768.639672845193
Rh001_041_013+    i_041    tia_h_in_001_013+    15164.652563252863
Rh001_041_013-    i_041    tia_h_in_001_013-    13891.234851748295
Rh001_042_013+    i_042    tia_h_in_001_013+    14338.30910309509
Rh001_042_013-    i_042    tia_h_in_001_013-    14864.945161425741
Rh001_043_013+    i_043    tia_h_in_001_013+    15184.066745613394
Rh001_043_013-    i_043    tia_h_in_001_013-    15115.204628807565
Rh001_044_013+    i_044    tia_h_in_001_013+    14749.15543334519
Rh001_044_013-    i_044    tia_h_in_001_013-    14966.608459738563
Rh001_045_013+    i_045    tia_h_in_001_013+    11871.22601317317
Rh001_045_013-    i_045    tia_h_in_001_013-    15197.141718913503
Rh001_046_013+    i_046    tia_h_in_001_013+    12205.4944258556
Rh001_046_013-    i_046    tia_h_in_001_013-    15000
Rh001_047_013+    i_047    tia_h_in_001_013+    15000
Rh001_047_013-    i_047    tia_h_in_001_013-    14893.868222636736
Rh001_048_013+    i_048    tia_h_in_001_013+    14784.905901747532
Rh001_048_013-    i_048    tia_h_in_001_013-    14533.990143086077
Rh001_049_013+    i_049    tia_h_in_001_013+    14980.662660142047
Rh001_049_013-    i_049    tia_h_in_001_013-    13956.53404364807
Rh001_050_013+    i_050    tia_h_in_001_013+    14961.887542683295
Rh001_050_013-    i_050    tia_h_in_001_013-    14879.201623905754
Rh001_051_013+    i_051    tia_h_in_001_013+    14796.74916156922
Rh001_051_013-    i_051    tia_h_in_001_013-    15135.792573816634
Rh001_052_013+    i_052    tia_h_in_001_013+    14775.987879987006
Rh001_052_013-    i_052    tia_h_in_001_013-    13546.616232320928
Rh001_053_013+    i_053    tia_h_in_001_013+    14836.532646825111
Rh001_053_013-    i_053    tia_h_in_001_013-    13603.447764368346
Rh001_054_013+    i_054    tia_h_in_001_013+    13645.344810686847
Rh001_054_013-    i_054    tia_h_in_001_013-    14870.788615060274
Rh001_055_013+    i_055    tia_h_in_001_013+    14013.817946976176
Rh001_055_013-    i_055    tia_h_in_001_013-    15025.55169507553
Rh001_056_013+    i_056    tia_h_in_001_013+    14718.689264190061
Rh001_056_013-    i_056    tia_h_in_001_013-    15098.558995549694
Rh001_057_013+    i_057    tia_h_in_001_013+    15000
Rh001_057_013-    i_057    tia_h_in_001_013-    14935.389060154785
Rh001_058_013+    i_058    tia_h_in_001_013+    14974.473933623487
Rh001_058_013-    i_058    tia_h_in_001_013-    14205.535122710988
Rh001_059_013+    i_059    tia_h_in_001_013+    14892.622353057055
Rh001_059_013-    i_059    tia_h_in_001_013-    14375.107073669395
Rh001_060_013+    i_060    tia_h_in_001_013+    15000
Rh001_060_013-    i_060    tia_h_in_001_013-    15195.270995328168
Rh001_061_013+    i_061    tia_h_in_001_013+    14941.468401524024
Rh001_061_013-    i_061    tia_h_in_001_013-    14640.97124609266
Rh001_062_013+    i_062    tia_h_in_001_013+    14796.786748498524
Rh001_062_013-    i_062    tia_h_in_001_013-    14336.198640406355
Rh001_063_013+    i_063    tia_h_in_001_013+    15064.813822418153
Rh001_063_013-    i_063    tia_h_in_001_013-    13268.847097365417
Rh001_064_013+    i_064    tia_h_in_001_013+    13274.865062403405
Rh001_064_013-    i_064    tia_h_in_001_013-    15000

* Neuron 14
Rh001_001_014+    i_001    tia_h_in_001_014+    15082.176599406173
Rh001_001_014-    i_001    tia_h_in_001_014-    13827.583237232566
Rh001_002_014+    i_002    tia_h_in_001_014+    15046.190849265779
Rh001_002_014-    i_002    tia_h_in_001_014-    14491.372385809012
Rh001_003_014+    i_003    tia_h_in_001_014+    14891.666708676255
Rh001_003_014-    i_003    tia_h_in_001_014-    14927.082088054469
Rh001_004_014+    i_004    tia_h_in_001_014+    14952.107264081806
Rh001_004_014-    i_004    tia_h_in_001_014-    14049.635134329672
Rh001_005_014+    i_005    tia_h_in_001_014+    5000
Rh001_005_014-    i_005    tia_h_in_001_014-    15085.106175577224
Rh001_006_014+    i_006    tia_h_in_001_014+    14848.48207865927
Rh001_006_014-    i_006    tia_h_in_001_014-    13120.929524530698
Rh001_007_014+    i_007    tia_h_in_001_014+    15100.897103300078
Rh001_007_014-    i_007    tia_h_in_001_014-    13698.254106223316
Rh001_008_014+    i_008    tia_h_in_001_014+    5000
Rh001_008_014-    i_008    tia_h_in_001_014-    13457.92769359438
Rh001_009_014+    i_009    tia_h_in_001_014+    15046.792667406839
Rh001_009_014-    i_009    tia_h_in_001_014-    14301.212088135851
Rh001_010_014+    i_010    tia_h_in_001_014+    15192.334978209728
Rh001_010_014-    i_010    tia_h_in_001_014-    14198.872660369232
Rh001_011_014+    i_011    tia_h_in_001_014+    15155.056309020216
Rh001_011_014-    i_011    tia_h_in_001_014-    15049.507265075626
Rh001_012_014+    i_012    tia_h_in_001_014+    15021.848877522285
Rh001_012_014-    i_012    tia_h_in_001_014-    14449.980729767545
Rh001_013_014+    i_013    tia_h_in_001_014+    14429.170850357184
Rh001_013_014-    i_013    tia_h_in_001_014-    14834.26205564966
Rh001_014_014+    i_014    tia_h_in_001_014+    13900.285236559448
Rh001_014_014-    i_014    tia_h_in_001_014-    5000
Rh001_015_014+    i_015    tia_h_in_001_014+    14875.602504594302
Rh001_015_014-    i_015    tia_h_in_001_014-    14838.138974723946
Rh001_016_014+    i_016    tia_h_in_001_014+    14709.440132975482
Rh001_016_014-    i_016    tia_h_in_001_014-    13937.946429178199
Rh001_017_014+    i_017    tia_h_in_001_014+    15123.753109000078
Rh001_017_014-    i_017    tia_h_in_001_014-    13494.404979110845
Rh001_018_014+    i_018    tia_h_in_001_014+    14510.915525010942
Rh001_018_014-    i_018    tia_h_in_001_014-    15052.545884780184
Rh001_019_014+    i_019    tia_h_in_001_014+    14993.561744419547
Rh001_019_014-    i_019    tia_h_in_001_014-    14249.978704965488
Rh001_020_014+    i_020    tia_h_in_001_014+    5000
Rh001_020_014-    i_020    tia_h_in_001_014-    14955.94413283347
Rh001_021_014+    i_021    tia_h_in_001_014+    14284.674669761876
Rh001_021_014-    i_021    tia_h_in_001_014-    14894.24015710085
Rh001_022_014+    i_022    tia_h_in_001_014+    14720.222353431256
Rh001_022_014-    i_022    tia_h_in_001_014-    15035.989274141568
Rh001_023_014+    i_023    tia_h_in_001_014+    13928.998518485847
Rh001_023_014-    i_023    tia_h_in_001_014-    14875.255567423594
Rh001_024_014+    i_024    tia_h_in_001_014+    13896.19088529462
Rh001_024_014-    i_024    tia_h_in_001_014-    15194.48784020063
Rh001_025_014+    i_025    tia_h_in_001_014+    14948.643100011708
Rh001_025_014-    i_025    tia_h_in_001_014-    15089.631833777681
Rh001_026_014+    i_026    tia_h_in_001_014+    15108.193585315588
Rh001_026_014-    i_026    tia_h_in_001_014-    13604.111961692044
Rh001_027_014+    i_027    tia_h_in_001_014+    15000
Rh001_027_014-    i_027    tia_h_in_001_014-    15175.589126163213
Rh001_028_014+    i_028    tia_h_in_001_014+    14870.904716454535
Rh001_028_014-    i_028    tia_h_in_001_014-    15000
Rh001_029_014+    i_029    tia_h_in_001_014+    15131.109473293527
Rh001_029_014-    i_029    tia_h_in_001_014-    13864.123979172811
Rh001_030_014+    i_030    tia_h_in_001_014+    14148.585091762243
Rh001_030_014-    i_030    tia_h_in_001_014-    14992.334069191644
Rh001_031_014+    i_031    tia_h_in_001_014+    14029.482046934037
Rh001_031_014-    i_031    tia_h_in_001_014-    15147.554484101369
Rh001_032_014+    i_032    tia_h_in_001_014+    15090.248869099156
Rh001_032_014-    i_032    tia_h_in_001_014-    14940.51142297736
Rh001_033_014+    i_033    tia_h_in_001_014+    15013.79638869361
Rh001_033_014-    i_033    tia_h_in_001_014-    14627.571823933571
Rh001_034_014+    i_034    tia_h_in_001_014+    15033.559181514729
Rh001_034_014-    i_034    tia_h_in_001_014-    13680.927607784688
Rh001_035_014+    i_035    tia_h_in_001_014+    15024.488016166883
Rh001_035_014-    i_035    tia_h_in_001_014-    14665.597533112692
Rh001_036_014+    i_036    tia_h_in_001_014+    13548.225187463875
Rh001_036_014-    i_036    tia_h_in_001_014-    5000
Rh001_037_014+    i_037    tia_h_in_001_014+    14702.498353949542
Rh001_037_014-    i_037    tia_h_in_001_014-    14982.394020880649
Rh001_038_014+    i_038    tia_h_in_001_014+    15024.81443020917
Rh001_038_014-    i_038    tia_h_in_001_014-    14965.705469539964
Rh001_039_014+    i_039    tia_h_in_001_014+    5000
Rh001_039_014-    i_039    tia_h_in_001_014-    14386.002129302704
Rh001_040_014+    i_040    tia_h_in_001_014+    15048.18492369162
Rh001_040_014-    i_040    tia_h_in_001_014-    14195.845325938164
Rh001_041_014+    i_041    tia_h_in_001_014+    14519.878152047479
Rh001_041_014-    i_041    tia_h_in_001_014-    14984.842125772246
Rh001_042_014+    i_042    tia_h_in_001_014+    15067.949066664818
Rh001_042_014-    i_042    tia_h_in_001_014-    14613.255629428026
Rh001_043_014+    i_043    tia_h_in_001_014+    14256.05176275704
Rh001_043_014-    i_043    tia_h_in_001_014-    14982.055002256422
Rh001_044_014+    i_044    tia_h_in_001_014+    15066.61893011208
Rh001_044_014-    i_044    tia_h_in_001_014-    14621.961246524246
Rh001_045_014+    i_045    tia_h_in_001_014+    14656.349448054245
Rh001_045_014-    i_045    tia_h_in_001_014-    14968.462553742038
Rh001_046_014+    i_046    tia_h_in_001_014+    14719.475537406293
Rh001_046_014-    i_046    tia_h_in_001_014-    14978.251922368272
Rh001_047_014+    i_047    tia_h_in_001_014+    15089.77045680287
Rh001_047_014-    i_047    tia_h_in_001_014-    15130.058831983071
Rh001_048_014+    i_048    tia_h_in_001_014+    15000
Rh001_048_014-    i_048    tia_h_in_001_014-    15000
Rh001_049_014+    i_049    tia_h_in_001_014+    14427.447467758631
Rh001_049_014-    i_049    tia_h_in_001_014-    15042.368244378431
Rh001_050_014+    i_050    tia_h_in_001_014+    13953.701097580784
Rh001_050_014-    i_050    tia_h_in_001_014-    14793.01282637236
Rh001_051_014+    i_051    tia_h_in_001_014+    14178.01106130479
Rh001_051_014-    i_051    tia_h_in_001_014-    5000
Rh001_052_014+    i_052    tia_h_in_001_014+    14908.334211947484
Rh001_052_014-    i_052    tia_h_in_001_014-    14322.180614271256
Rh001_053_014+    i_053    tia_h_in_001_014+    15019.414739972237
Rh001_053_014-    i_053    tia_h_in_001_014-    13477.527033554874
Rh001_054_014+    i_054    tia_h_in_001_014+    5000
Rh001_054_014-    i_054    tia_h_in_001_014-    14998.71507470208
Rh001_055_014+    i_055    tia_h_in_001_014+    5000
Rh001_055_014-    i_055    tia_h_in_001_014-    14820.479225037841
Rh001_056_014+    i_056    tia_h_in_001_014+    14993.416674742133
Rh001_056_014-    i_056    tia_h_in_001_014-    14404.461724388453
Rh001_057_014+    i_057    tia_h_in_001_014+    15113.388690929407
Rh001_057_014-    i_057    tia_h_in_001_014-    14357.737596276207
Rh001_058_014+    i_058    tia_h_in_001_014+    15146.961153117929
Rh001_058_014-    i_058    tia_h_in_001_014-    14480.819223980103
Rh001_059_014+    i_059    tia_h_in_001_014+    14016.025430666068
Rh001_059_014-    i_059    tia_h_in_001_014-    14961.274060002183
Rh001_060_014+    i_060    tia_h_in_001_014+    15130.925973832784
Rh001_060_014-    i_060    tia_h_in_001_014-    15238.05649887246
Rh001_061_014+    i_061    tia_h_in_001_014+    15095.249674227525
Rh001_061_014-    i_061    tia_h_in_001_014-    14168.973493802703
Rh001_062_014+    i_062    tia_h_in_001_014+    15013.050672824254
Rh001_062_014-    i_062    tia_h_in_001_014-    14202.337288566892
Rh001_063_014+    i_063    tia_h_in_001_014+    14965.271397910808
Rh001_063_014-    i_063    tia_h_in_001_014-    14488.28585285205
Rh001_064_014+    i_064    tia_h_in_001_014+    14993.76749730229
Rh001_064_014-    i_064    tia_h_in_001_014-    14123.995736254068

* Neuron 15
Rh001_001_015+    i_001    tia_h_in_001_015+    13619.416178476738
Rh001_001_015-    i_001    tia_h_in_001_015-    5000
Rh001_002_015+    i_002    tia_h_in_001_015+    14321.7536141874
Rh001_002_015-    i_002    tia_h_in_001_015-    15002.168382093741
Rh001_003_015+    i_003    tia_h_in_001_015+    13866.414545244814
Rh001_003_015-    i_003    tia_h_in_001_015-    14906.589117522903
Rh001_004_015+    i_004    tia_h_in_001_015+    15044.534832858426
Rh001_004_015-    i_004    tia_h_in_001_015-    14891.038769322395
Rh001_005_015+    i_005    tia_h_in_001_015+    14997.339499443568
Rh001_005_015-    i_005    tia_h_in_001_015-    15194.891756105771
Rh001_006_015+    i_006    tia_h_in_001_015+    15000
Rh001_006_015-    i_006    tia_h_in_001_015-    14946.850511953393
Rh001_007_015+    i_007    tia_h_in_001_015+    14980.131892102481
Rh001_007_015-    i_007    tia_h_in_001_015-    13575.334780901407
Rh001_008_015+    i_008    tia_h_in_001_015+    15275.861203191918
Rh001_008_015-    i_008    tia_h_in_001_015-    14907.321938896283
Rh001_009_015+    i_009    tia_h_in_001_015+    14995.554316247077
Rh001_009_015-    i_009    tia_h_in_001_015-    14758.634778023521
Rh001_010_015+    i_010    tia_h_in_001_015+    15000
Rh001_010_015-    i_010    tia_h_in_001_015-    13909.639721487103
Rh001_011_015+    i_011    tia_h_in_001_015+    15027.521684995996
Rh001_011_015-    i_011    tia_h_in_001_015-    13745.528023486879
Rh001_012_015+    i_012    tia_h_in_001_015+    13932.27275566141
Rh001_012_015-    i_012    tia_h_in_001_015-    15047.125866053388
Rh001_013_015+    i_013    tia_h_in_001_015+    13981.608542842614
Rh001_013_015-    i_013    tia_h_in_001_015-    14875.736895188727
Rh001_014_015+    i_014    tia_h_in_001_015+    14448.893475432365
Rh001_014_015-    i_014    tia_h_in_001_015-    14928.601799399088
Rh001_015_015+    i_015    tia_h_in_001_015+    13812.316553905039
Rh001_015_015-    i_015    tia_h_in_001_015-    15025.939847200121
Rh001_016_015+    i_016    tia_h_in_001_015+    14944.568345432728
Rh001_016_015-    i_016    tia_h_in_001_015-    14400.459446381014
Rh001_017_015+    i_017    tia_h_in_001_015+    14964.567381143695
Rh001_017_015-    i_017    tia_h_in_001_015-    14747.645204265245
Rh001_018_015+    i_018    tia_h_in_001_015+    14628.062121707742
Rh001_018_015-    i_018    tia_h_in_001_015-    14909.334202570082
Rh001_019_015+    i_019    tia_h_in_001_015+    14833.766125054528
Rh001_019_015-    i_019    tia_h_in_001_015-    14806.16380713591
Rh001_020_015+    i_020    tia_h_in_001_015+    15147.313518569978
Rh001_020_015-    i_020    tia_h_in_001_015-    5000
Rh001_021_015+    i_021    tia_h_in_001_015+    5000
Rh001_021_015-    i_021    tia_h_in_001_015-    13650.418591630774
Rh001_022_015+    i_022    tia_h_in_001_015+    14938.357537711887
Rh001_022_015-    i_022    tia_h_in_001_015-    15135.422992443908
Rh001_023_015+    i_023    tia_h_in_001_015+    15035.391880540268
Rh001_023_015-    i_023    tia_h_in_001_015-    13908.212301439491
Rh001_024_015+    i_024    tia_h_in_001_015+    5000
Rh001_024_015-    i_024    tia_h_in_001_015-    15034.744526056988
Rh001_025_015+    i_025    tia_h_in_001_015+    13641.734849562783
Rh001_025_015-    i_025    tia_h_in_001_015-    15103.930496936066
Rh001_026_015+    i_026    tia_h_in_001_015+    5000
Rh001_026_015-    i_026    tia_h_in_001_015-    14335.655080077157
Rh001_027_015+    i_027    tia_h_in_001_015+    15108.079501340073
Rh001_027_015-    i_027    tia_h_in_001_015-    14486.695939909434
Rh001_028_015+    i_028    tia_h_in_001_015+    14243.972946326301
Rh001_028_015-    i_028    tia_h_in_001_015-    14912.872083805296
Rh001_029_015+    i_029    tia_h_in_001_015+    15267.66259237067
Rh001_029_015-    i_029    tia_h_in_001_015-    14176.151563640668
Rh001_030_015+    i_030    tia_h_in_001_015+    14908.934166589368
Rh001_030_015-    i_030    tia_h_in_001_015-    14710.106812576154
Rh001_031_015+    i_031    tia_h_in_001_015+    13778.034251421912
Rh001_031_015-    i_031    tia_h_in_001_015-    14987.872943956982
Rh001_032_015+    i_032    tia_h_in_001_015+    14759.437621070467
Rh001_032_015-    i_032    tia_h_in_001_015-    14359.661470377732
Rh001_033_015+    i_033    tia_h_in_001_015+    15073.059977022702
Rh001_033_015-    i_033    tia_h_in_001_015-    13969.347868846116
Rh001_034_015+    i_034    tia_h_in_001_015+    15079.560145839552
Rh001_034_015-    i_034    tia_h_in_001_015-    13960.546122671138
Rh001_035_015+    i_035    tia_h_in_001_015+    15010.93032124239
Rh001_035_015-    i_035    tia_h_in_001_015-    14615.514840498296
Rh001_036_015+    i_036    tia_h_in_001_015+    14975.731892760901
Rh001_036_015-    i_036    tia_h_in_001_015-    14082.714938234461
Rh001_037_015+    i_037    tia_h_in_001_015+    15159.61921792163
Rh001_037_015-    i_037    tia_h_in_001_015-    5000
Rh001_038_015+    i_038    tia_h_in_001_015+    14316.961834025637
Rh001_038_015-    i_038    tia_h_in_001_015-    15041.524914127649
Rh001_039_015+    i_039    tia_h_in_001_015+    14729.305572961883
Rh001_039_015-    i_039    tia_h_in_001_015-    15015.046628624392
Rh001_040_015+    i_040    tia_h_in_001_015+    15024.069723387664
Rh001_040_015-    i_040    tia_h_in_001_015-    14287.366539658131
Rh001_041_015+    i_041    tia_h_in_001_015+    15200.966876701317
Rh001_041_015-    i_041    tia_h_in_001_015-    13887.982131698785
Rh001_042_015+    i_042    tia_h_in_001_015+    15064.05852011654
Rh001_042_015-    i_042    tia_h_in_001_015-    14299.833327673341
Rh001_043_015+    i_043    tia_h_in_001_015+    15021.499269872165
Rh001_043_015-    i_043    tia_h_in_001_015-    14240.705171133726
Rh001_044_015+    i_044    tia_h_in_001_015+    14938.989217999504
Rh001_044_015-    i_044    tia_h_in_001_015-    14406.474341711888
Rh001_045_015+    i_045    tia_h_in_001_015+    14922.573347701655
Rh001_045_015-    i_045    tia_h_in_001_015-    13633.555176835252
Rh001_046_015+    i_046    tia_h_in_001_015+    14741.641084211331
Rh001_046_015-    i_046    tia_h_in_001_015-    14872.96669609111
Rh001_047_015+    i_047    tia_h_in_001_015+    14988.496371833258
Rh001_047_015-    i_047    tia_h_in_001_015-    14013.344044605154
Rh001_048_015+    i_048    tia_h_in_001_015+    15000
Rh001_048_015-    i_048    tia_h_in_001_015-    13596.506817849688
Rh001_049_015+    i_049    tia_h_in_001_015+    15133.487464406113
Rh001_049_015-    i_049    tia_h_in_001_015-    13664.795095651474
Rh001_050_015+    i_050    tia_h_in_001_015+    15000
Rh001_050_015-    i_050    tia_h_in_001_015-    15057.762700372392
Rh001_051_015+    i_051    tia_h_in_001_015+    14850.900365152123
Rh001_051_015-    i_051    tia_h_in_001_015-    14130.32867410991
Rh001_052_015+    i_052    tia_h_in_001_015+    15206.785367552033
Rh001_052_015-    i_052    tia_h_in_001_015-    14262.896350906945
Rh001_053_015+    i_053    tia_h_in_001_015+    14047.378135080438
Rh001_053_015-    i_053    tia_h_in_001_015-    15215.012195848114
Rh001_054_015+    i_054    tia_h_in_001_015+    14264.341820731534
Rh001_054_015-    i_054    tia_h_in_001_015-    14705.357954010175
Rh001_055_015+    i_055    tia_h_in_001_015+    14231.096423187364
Rh001_055_015-    i_055    tia_h_in_001_015-    15116.71482535034
Rh001_056_015+    i_056    tia_h_in_001_015+    15103.359642619023
Rh001_056_015-    i_056    tia_h_in_001_015-    13567.953315346122
Rh001_057_015+    i_057    tia_h_in_001_015+    5000
Rh001_057_015-    i_057    tia_h_in_001_015-    5000
Rh001_058_015+    i_058    tia_h_in_001_015+    14864.939922941132
Rh001_058_015-    i_058    tia_h_in_001_015-    14222.517959374274
Rh001_059_015+    i_059    tia_h_in_001_015+    14108.895903504565
Rh001_059_015-    i_059    tia_h_in_001_015-    15062.128602725918
Rh001_060_015+    i_060    tia_h_in_001_015+    14825.639786772927
Rh001_060_015-    i_060    tia_h_in_001_015-    14761.991262746677
Rh001_061_015+    i_061    tia_h_in_001_015+    14745.654767647999
Rh001_061_015-    i_061    tia_h_in_001_015-    13700.625357244693
Rh001_062_015+    i_062    tia_h_in_001_015+    5000
Rh001_062_015-    i_062    tia_h_in_001_015-    14912.581698697371
Rh001_063_015+    i_063    tia_h_in_001_015+    15000
Rh001_063_015-    i_063    tia_h_in_001_015-    13548.551321853527
Rh001_064_015+    i_064    tia_h_in_001_015+    15090.084021909763
Rh001_064_015-    i_064    tia_h_in_001_015-    14585.61206599066

* Neuron 16
Rh001_001_016+    i_001    tia_h_in_001_016+    11658.139884886765
Rh001_001_016-    i_001    tia_h_in_001_016-    14962.182208520946
Rh001_002_016+    i_002    tia_h_in_001_016+    11296.100014836145
Rh001_002_016-    i_002    tia_h_in_001_016-    15000
Rh001_003_016+    i_003    tia_h_in_001_016+    14311.022461121784
Rh001_003_016-    i_003    tia_h_in_001_016-    15101.904043381714
Rh001_004_016+    i_004    tia_h_in_001_016+    15000
Rh001_004_016-    i_004    tia_h_in_001_016-    13086.680103190592
Rh001_005_016+    i_005    tia_h_in_001_016+    15065.538671183635
Rh001_005_016-    i_005    tia_h_in_001_016-    10513.674114336316
Rh001_006_016+    i_006    tia_h_in_001_016+    15051.283328040561
Rh001_006_016-    i_006    tia_h_in_001_016-    9950.272675069025
Rh001_007_016+    i_007    tia_h_in_001_016+    14973.927872013262
Rh001_007_016-    i_007    tia_h_in_001_016-    14602.121730494224
Rh001_008_016+    i_008    tia_h_in_001_016+    5000
Rh001_008_016-    i_008    tia_h_in_001_016-    15070.741315637606
Rh001_009_016+    i_009    tia_h_in_001_016+    15044.77700122375
Rh001_009_016-    i_009    tia_h_in_001_016-    14115.521895426868
Rh001_010_016+    i_010    tia_h_in_001_016+    14944.351305963122
Rh001_010_016-    i_010    tia_h_in_001_016-    15000
Rh001_011_016+    i_011    tia_h_in_001_016+    15136.714640951985
Rh001_011_016-    i_011    tia_h_in_001_016-    13296.038395717575
Rh001_012_016+    i_012    tia_h_in_001_016+    15053.214200589451
Rh001_012_016-    i_012    tia_h_in_001_016-    13101.453155915773
Rh001_013_016+    i_013    tia_h_in_001_016+    14942.328433199116
Rh001_013_016-    i_013    tia_h_in_001_016-    14439.324971830289
Rh001_014_016+    i_014    tia_h_in_001_016+    14578.513100450431
Rh001_014_016-    i_014    tia_h_in_001_016-    15081.458455268235
Rh001_015_016+    i_015    tia_h_in_001_016+    15000
Rh001_015_016-    i_015    tia_h_in_001_016-    15042.157157410486
Rh001_016_016+    i_016    tia_h_in_001_016+    12810.491535261373
Rh001_016_016-    i_016    tia_h_in_001_016-    15146.149214887395
Rh001_017_016+    i_017    tia_h_in_001_016+    15194.281598998194
Rh001_017_016-    i_017    tia_h_in_001_016-    15018.79310976798
Rh001_018_016+    i_018    tia_h_in_001_016+    13089.360242349558
Rh001_018_016-    i_018    tia_h_in_001_016-    15000
Rh001_019_016+    i_019    tia_h_in_001_016+    14956.154339429973
Rh001_019_016-    i_019    tia_h_in_001_016-    14703.35909650228
Rh001_020_016+    i_020    tia_h_in_001_016+    5000
Rh001_020_016-    i_020    tia_h_in_001_016-    13391.828444740964
Rh001_021_016+    i_021    tia_h_in_001_016+    15055.34572064621
Rh001_021_016-    i_021    tia_h_in_001_016-    12337.957394075727
Rh001_022_016+    i_022    tia_h_in_001_016+    15173.383861210132
Rh001_022_016-    i_022    tia_h_in_001_016-    14853.369274774608
Rh001_023_016+    i_023    tia_h_in_001_016+    15107.74817985707
Rh001_023_016-    i_023    tia_h_in_001_016-    13715.603417809774
Rh001_024_016+    i_024    tia_h_in_001_016+    5000
Rh001_024_016-    i_024    tia_h_in_001_016-    15061.846298315542
Rh001_025_016+    i_025    tia_h_in_001_016+    5000
Rh001_025_016-    i_025    tia_h_in_001_016-    15082.452517723972
Rh001_026_016+    i_026    tia_h_in_001_016+    14941.876578165737
Rh001_026_016-    i_026    tia_h_in_001_016-    13981.327881301586
Rh001_027_016+    i_027    tia_h_in_001_016+    15172.93957740518
Rh001_027_016-    i_027    tia_h_in_001_016-    14023.723202268413
Rh001_028_016+    i_028    tia_h_in_001_016+    14931.380249578253
Rh001_028_016-    i_028    tia_h_in_001_016-    14450.210034771917
Rh001_029_016+    i_029    tia_h_in_001_016+    14913.87881151721
Rh001_029_016-    i_029    tia_h_in_001_016-    15032.011534610967
Rh001_030_016+    i_030    tia_h_in_001_016+    14938.526685451885
Rh001_030_016-    i_030    tia_h_in_001_016-    14572.198313153855
Rh001_031_016+    i_031    tia_h_in_001_016+    13251.586096432695
Rh001_031_016-    i_031    tia_h_in_001_016-    15096.287575994435
Rh001_032_016+    i_032    tia_h_in_001_016+    13670.488672290392
Rh001_032_016-    i_032    tia_h_in_001_016-    15071.480940639927
Rh001_033_016+    i_033    tia_h_in_001_016+    14963.840714558464
Rh001_033_016-    i_033    tia_h_in_001_016-    14817.138506838426
Rh001_034_016+    i_034    tia_h_in_001_016+    15034.310488649151
Rh001_034_016-    i_034    tia_h_in_001_016-    14882.55913079213
Rh001_035_016+    i_035    tia_h_in_001_016+    14970.121013376756
Rh001_035_016-    i_035    tia_h_in_001_016-    12950.422894944048
Rh001_036_016+    i_036    tia_h_in_001_016+    14917.196813791128
Rh001_036_016-    i_036    tia_h_in_001_016-    12597.28998651083
Rh001_037_016+    i_037    tia_h_in_001_016+    14228.819372698727
Rh001_037_016-    i_037    tia_h_in_001_016-    14948.514620354013
Rh001_038_016+    i_038    tia_h_in_001_016+    12543.244589573213
Rh001_038_016-    i_038    tia_h_in_001_016-    14965.131856879194
Rh001_039_016+    i_039    tia_h_in_001_016+    14410.153984956696
Rh001_039_016-    i_039    tia_h_in_001_016-    15025.26092621568
Rh001_040_016+    i_040    tia_h_in_001_016+    13001.5697920221
Rh001_040_016-    i_040    tia_h_in_001_016-    15011.478024988819
Rh001_041_016+    i_041    tia_h_in_001_016+    15107.28845053291
Rh001_041_016-    i_041    tia_h_in_001_016-    13044.387238537794
Rh001_042_016+    i_042    tia_h_in_001_016+    14997.181602691848
Rh001_042_016-    i_042    tia_h_in_001_016-    13851.722259029732
Rh001_043_016+    i_043    tia_h_in_001_016+    14971.746041361635
Rh001_043_016-    i_043    tia_h_in_001_016-    5000
Rh001_044_016+    i_044    tia_h_in_001_016+    12691.92177131071
Rh001_044_016-    i_044    tia_h_in_001_016-    14847.410836035002
Rh001_045_016+    i_045    tia_h_in_001_016+    12624.481147232422
Rh001_045_016-    i_045    tia_h_in_001_016-    15141.024043814714
Rh001_046_016+    i_046    tia_h_in_001_016+    12961.121434896631
Rh001_046_016-    i_046    tia_h_in_001_016-    14852.884341582589
Rh001_047_016+    i_047    tia_h_in_001_016+    14049.09020709615
Rh001_047_016-    i_047    tia_h_in_001_016-    14818.447361799379
Rh001_048_016+    i_048    tia_h_in_001_016+    14846.767238019593
Rh001_048_016-    i_048    tia_h_in_001_016-    12833.415447145337
Rh001_049_016+    i_049    tia_h_in_001_016+    15000
Rh001_049_016-    i_049    tia_h_in_001_016-    5000
Rh001_050_016+    i_050    tia_h_in_001_016+    14980.527867022194
Rh001_050_016-    i_050    tia_h_in_001_016-    12879.723475659774
Rh001_051_016+    i_051    tia_h_in_001_016+    15188.009173109394
Rh001_051_016-    i_051    tia_h_in_001_016-    13234.52508626637
Rh001_052_016+    i_052    tia_h_in_001_016+    13762.683909996273
Rh001_052_016-    i_052    tia_h_in_001_016-    14951.651497282419
Rh001_053_016+    i_053    tia_h_in_001_016+    13381.520545261754
Rh001_053_016-    i_053    tia_h_in_001_016-    15024.191380305334
Rh001_054_016+    i_054    tia_h_in_001_016+    12010.384928193129
Rh001_054_016-    i_054    tia_h_in_001_016-    14839.789630050474
Rh001_055_016+    i_055    tia_h_in_001_016+    13442.633170788637
Rh001_055_016-    i_055    tia_h_in_001_016-    15000
Rh001_056_016+    i_056    tia_h_in_001_016+    15032.146369512759
Rh001_056_016-    i_056    tia_h_in_001_016-    13828.84996558483
Rh001_057_016+    i_057    tia_h_in_001_016+    15157.252526447397
Rh001_057_016-    i_057    tia_h_in_001_016-    12819.843243325617
Rh001_058_016+    i_058    tia_h_in_001_016+    14950.560433765808
Rh001_058_016-    i_058    tia_h_in_001_016-    14025.027022425578
Rh001_059_016+    i_059    tia_h_in_001_016+    11629.17495058309
Rh001_059_016-    i_059    tia_h_in_001_016-    15000
Rh001_060_016+    i_060    tia_h_in_001_016+    10931.720969956272
Rh001_060_016-    i_060    tia_h_in_001_016-    14967.087363700526
Rh001_061_016+    i_061    tia_h_in_001_016+    11324.545652543802
Rh001_061_016-    i_061    tia_h_in_001_016-    15096.17170752916
Rh001_062_016+    i_062    tia_h_in_001_016+    15065.70416188977
Rh001_062_016-    i_062    tia_h_in_001_016-    14722.58986393884
Rh001_063_016+    i_063    tia_h_in_001_016+    15028.241776087305
Rh001_063_016-    i_063    tia_h_in_001_016-    11394.300164833392
Rh001_064_016+    i_064    tia_h_in_001_016+    15000
Rh001_064_016-    i_064    tia_h_in_001_016-    11291.382964900347

* Neuron 17
Rh001_001_017+    i_001    tia_h_in_001_017+    14849.366840252795
Rh001_001_017-    i_001    tia_h_in_001_017-    13233.205143990737
Rh001_002_017+    i_002    tia_h_in_001_017+    14280.161541013595
Rh001_002_017-    i_002    tia_h_in_001_017-    14919.270162745152
Rh001_003_017+    i_003    tia_h_in_001_017+    15033.407305748458
Rh001_003_017-    i_003    tia_h_in_001_017-    11831.326180194503
Rh001_004_017+    i_004    tia_h_in_001_017+    14956.867809427344
Rh001_004_017-    i_004    tia_h_in_001_017-    8913.056258542869
Rh001_005_017+    i_005    tia_h_in_001_017+    15042.789768890894
Rh001_005_017-    i_005    tia_h_in_001_017-    15000
Rh001_006_017+    i_006    tia_h_in_001_017+    12549.238077086276
Rh001_006_017-    i_006    tia_h_in_001_017-    15011.726798337511
Rh001_007_017+    i_007    tia_h_in_001_017+    12053.503724583985
Rh001_007_017-    i_007    tia_h_in_001_017-    15000
Rh001_008_017+    i_008    tia_h_in_001_017+    12083.920235358892
Rh001_008_017-    i_008    tia_h_in_001_017-    15048.936228173816
Rh001_009_017+    i_009    tia_h_in_001_017+    15158.49021939782
Rh001_009_017-    i_009    tia_h_in_001_017-    14235.81942484671
Rh001_010_017+    i_010    tia_h_in_001_017+    14788.916008395638
Rh001_010_017-    i_010    tia_h_in_001_017-    12751.544507670238
Rh001_011_017+    i_011    tia_h_in_001_017+    14985.76506955514
Rh001_011_017-    i_011    tia_h_in_001_017-    5000
Rh001_012_017+    i_012    tia_h_in_001_017+    14825.553946911183
Rh001_012_017-    i_012    tia_h_in_001_017-    13411.076333809757
Rh001_013_017+    i_013    tia_h_in_001_017+    13655.118110862226
Rh001_013_017-    i_013    tia_h_in_001_017-    15071.39142385493
Rh001_014_017+    i_014    tia_h_in_001_017+    11023.565680408869
Rh001_014_017-    i_014    tia_h_in_001_017-    14957.761053795006
Rh001_015_017+    i_015    tia_h_in_001_017+    14227.604099891347
Rh001_015_017-    i_015    tia_h_in_001_017-    14857.049700036918
Rh001_016_017+    i_016    tia_h_in_001_017+    14910.024573369941
Rh001_016_017-    i_016    tia_h_in_001_017-    14616.342608486113
Rh001_017_017+    i_017    tia_h_in_001_017+    14896.486600450997
Rh001_017_017-    i_017    tia_h_in_001_017-    14424.854197383323
Rh001_018_017+    i_018    tia_h_in_001_017+    14929.42145714815
Rh001_018_017-    i_018    tia_h_in_001_017-    5000
Rh001_019_017+    i_019    tia_h_in_001_017+    15148.404232472165
Rh001_019_017-    i_019    tia_h_in_001_017-    12293.8545563228
Rh001_020_017+    i_020    tia_h_in_001_017+    15078.938114824457
Rh001_020_017-    i_020    tia_h_in_001_017-    14645.550345875117
Rh001_021_017+    i_021    tia_h_in_001_017+    13007.228319883629
Rh001_021_017-    i_021    tia_h_in_001_017-    15054.779131499527
Rh001_022_017+    i_022    tia_h_in_001_017+    13812.184207698452
Rh001_022_017-    i_022    tia_h_in_001_017-    14873.888206910422
Rh001_023_017+    i_023    tia_h_in_001_017+    13412.745883657592
Rh001_023_017-    i_023    tia_h_in_001_017-    15223.999027457832
Rh001_024_017+    i_024    tia_h_in_001_017+    14898.074342828231
Rh001_024_017-    i_024    tia_h_in_001_017-    13495.838237730306
Rh001_025_017+    i_025    tia_h_in_001_017+    14374.654100539985
Rh001_025_017-    i_025    tia_h_in_001_017-    15000
Rh001_026_017+    i_026    tia_h_in_001_017+    14285.523149004335
Rh001_026_017-    i_026    tia_h_in_001_017-    14935.891218539424
Rh001_027_017+    i_027    tia_h_in_001_017+    13523.802387316498
Rh001_027_017-    i_027    tia_h_in_001_017-    15143.73822661407
Rh001_028_017+    i_028    tia_h_in_001_017+    11951.656002442056
Rh001_028_017-    i_028    tia_h_in_001_017-    14977.140278636878
Rh001_029_017+    i_029    tia_h_in_001_017+    10326.22335377706
Rh001_029_017-    i_029    tia_h_in_001_017-    15138.099241832479
Rh001_030_017+    i_030    tia_h_in_001_017+    12739.915304194197
Rh001_030_017-    i_030    tia_h_in_001_017-    15102.66891943833
Rh001_031_017+    i_031    tia_h_in_001_017+    15047.156341645554
Rh001_031_017-    i_031    tia_h_in_001_017-    11869.252232857254
Rh001_032_017+    i_032    tia_h_in_001_017+    15073.516044684293
Rh001_032_017-    i_032    tia_h_in_001_017-    13919.480002005608
Rh001_033_017+    i_033    tia_h_in_001_017+    14911.693057339033
Rh001_033_017-    i_033    tia_h_in_001_017-    14127.670081728334
Rh001_034_017+    i_034    tia_h_in_001_017+    14816.307591041481
Rh001_034_017-    i_034    tia_h_in_001_017-    11668.746350772506
Rh001_035_017+    i_035    tia_h_in_001_017+    11685.073573614458
Rh001_035_017-    i_035    tia_h_in_001_017-    14990.416060419022
Rh001_036_017+    i_036    tia_h_in_001_017+    10703.832859887896
Rh001_036_017-    i_036    tia_h_in_001_017-    15210.928823958478
Rh001_037_017+    i_037    tia_h_in_001_017+    5000
Rh001_037_017-    i_037    tia_h_in_001_017-    15023.955876910095
Rh001_038_017+    i_038    tia_h_in_001_017+    14167.049177337198
Rh001_038_017-    i_038    tia_h_in_001_017-    14950.782716895174
Rh001_039_017+    i_039    tia_h_in_001_017+    14998.91973807079
Rh001_039_017-    i_039    tia_h_in_001_017-    14225.726507463763
Rh001_040_017+    i_040    tia_h_in_001_017+    13718.372798693954
Rh001_040_017-    i_040    tia_h_in_001_017-    15000
Rh001_041_017+    i_041    tia_h_in_001_017+    14038.402164926576
Rh001_041_017-    i_041    tia_h_in_001_017-    15017.067132019392
Rh001_042_017+    i_042    tia_h_in_001_017+    13400.739537572494
Rh001_042_017-    i_042    tia_h_in_001_017-    14956.540976877457
Rh001_043_017+    i_043    tia_h_in_001_017+    5000
Rh001_043_017-    i_043    tia_h_in_001_017-    14809.114729301247
Rh001_044_017+    i_044    tia_h_in_001_017+    14191.761708817776
Rh001_044_017-    i_044    tia_h_in_001_017-    15000
Rh001_045_017+    i_045    tia_h_in_001_017+    15065.807888725805
Rh001_045_017-    i_045    tia_h_in_001_017-    15000
Rh001_046_017+    i_046    tia_h_in_001_017+    14928.993266558464
Rh001_046_017-    i_046    tia_h_in_001_017-    15000
Rh001_047_017+    i_047    tia_h_in_001_017+    14738.264026078548
Rh001_047_017-    i_047    tia_h_in_001_017-    14091.186107432912
Rh001_048_017+    i_048    tia_h_in_001_017+    15033.325819362579
Rh001_048_017-    i_048    tia_h_in_001_017-    14830.4591670883
Rh001_049_017+    i_049    tia_h_in_001_017+    14922.512798861992
Rh001_049_017-    i_049    tia_h_in_001_017-    13631.896421515916
Rh001_050_017+    i_050    tia_h_in_001_017+    5000
Rh001_050_017-    i_050    tia_h_in_001_017-    14892.45243153114
Rh001_051_017+    i_051    tia_h_in_001_017+    12802.01422751418
Rh001_051_017-    i_051    tia_h_in_001_017-    15000
Rh001_052_017+    i_052    tia_h_in_001_017+    13040.809767330567
Rh001_052_017-    i_052    tia_h_in_001_017-    14839.596347190978
Rh001_053_017+    i_053    tia_h_in_001_017+    14921.369725271052
Rh001_053_017-    i_053    tia_h_in_001_017-    14150.433244184
Rh001_054_017+    i_054    tia_h_in_001_017+    15008.598222699964
Rh001_054_017-    i_054    tia_h_in_001_017-    11520.656939198296
Rh001_055_017+    i_055    tia_h_in_001_017+    15090.104905168117
Rh001_055_017-    i_055    tia_h_in_001_017-    13473.880241118675
Rh001_056_017+    i_056    tia_h_in_001_017+    15081.704739354318
Rh001_056_017-    i_056    tia_h_in_001_017-    12745.709362861133
Rh001_057_017+    i_057    tia_h_in_001_017+    12940.839163325654
Rh001_057_017-    i_057    tia_h_in_001_017-    14796.025549210475
Rh001_058_017+    i_058    tia_h_in_001_017+    12073.324028838762
Rh001_058_017-    i_058    tia_h_in_001_017-    14927.148774102969
Rh001_059_017+    i_059    tia_h_in_001_017+    12294.207659532882
Rh001_059_017-    i_059    tia_h_in_001_017-    5000
Rh001_060_017+    i_060    tia_h_in_001_017+    15232.890577133729
Rh001_060_017-    i_060    tia_h_in_001_017-    12117.05747981223
Rh001_061_017+    i_061    tia_h_in_001_017+    14812.240197940762
Rh001_061_017-    i_061    tia_h_in_001_017-    9173.590159439429
Rh001_062_017+    i_062    tia_h_in_001_017+    15049.082077012048
Rh001_062_017-    i_062    tia_h_in_001_017-    12156.658967010473
Rh001_063_017+    i_063    tia_h_in_001_017+    13832.651627527022
Rh001_063_017-    i_063    tia_h_in_001_017-    14945.065002398575
Rh001_064_017+    i_064    tia_h_in_001_017+    14695.803349940683
Rh001_064_017-    i_064    tia_h_in_001_017-    14941.832653954836

* Neuron 18
Rh001_001_018+    i_001    tia_h_in_001_018+    14908.324036362039
Rh001_001_018-    i_001    tia_h_in_001_018-    12042.10212276785
Rh001_002_018+    i_002    tia_h_in_001_018+    15070.398674317516
Rh001_002_018-    i_002    tia_h_in_001_018-    11799.928811911954
Rh001_003_018+    i_003    tia_h_in_001_018+    14951.417444938495
Rh001_003_018-    i_003    tia_h_in_001_018-    14296.979364378107
Rh001_004_018+    i_004    tia_h_in_001_018+    14916.50202061587
Rh001_004_018-    i_004    tia_h_in_001_018-    15000
Rh001_005_018+    i_005    tia_h_in_001_018+    14736.889111121307
Rh001_005_018-    i_005    tia_h_in_001_018-    15209.222681386878
Rh001_006_018+    i_006    tia_h_in_001_018+    15056.722532874137
Rh001_006_018-    i_006    tia_h_in_001_018-    13914.866415838074
Rh001_007_018+    i_007    tia_h_in_001_018+    14485.621212734704
Rh001_007_018-    i_007    tia_h_in_001_018-    15010.422033298228
Rh001_008_018+    i_008    tia_h_in_001_018+    13713.293369720723
Rh001_008_018-    i_008    tia_h_in_001_018-    15000
Rh001_009_018+    i_009    tia_h_in_001_018+    15059.837963317943
Rh001_009_018-    i_009    tia_h_in_001_018-    12454.878627206013
Rh001_010_018+    i_010    tia_h_in_001_018+    14979.260060243463
Rh001_010_018-    i_010    tia_h_in_001_018-    5000
Rh001_011_018+    i_011    tia_h_in_001_018+    13804.415161188788
Rh001_011_018-    i_011    tia_h_in_001_018-    15000
Rh001_012_018+    i_012    tia_h_in_001_018+    13921.20446232409
Rh001_012_018-    i_012    tia_h_in_001_018-    15052.520052456934
Rh001_013_018+    i_013    tia_h_in_001_018+    5000
Rh001_013_018-    i_013    tia_h_in_001_018-    14838.73157112581
Rh001_014_018+    i_014    tia_h_in_001_018+    13535.543193766525
Rh001_014_018-    i_014    tia_h_in_001_018-    14889.31889289435
Rh001_015_018+    i_015    tia_h_in_001_018+    14135.208877421506
Rh001_015_018-    i_015    tia_h_in_001_018-    14941.680082010967
Rh001_016_018+    i_016    tia_h_in_001_018+    14698.000994242997
Rh001_016_018-    i_016    tia_h_in_001_018-    13236.354303770551
Rh001_017_018+    i_017    tia_h_in_001_018+    14643.052849950249
Rh001_017_018-    i_017    tia_h_in_001_018-    14785.18143755838
Rh001_018_018+    i_018    tia_h_in_001_018+    14428.09920844195
Rh001_018_018-    i_018    tia_h_in_001_018-    15042.741830097393
Rh001_019_018+    i_019    tia_h_in_001_018+    5000
Rh001_019_018-    i_019    tia_h_in_001_018-    15097.951007099855
Rh001_020_018+    i_020    tia_h_in_001_018+    15190.765434764402
Rh001_020_018-    i_020    tia_h_in_001_018-    13970.49685040053
Rh001_021_018+    i_021    tia_h_in_001_018+    14303.55747189357
Rh001_021_018-    i_021    tia_h_in_001_018-    15301.965429830147
Rh001_022_018+    i_022    tia_h_in_001_018+    15014.83681433602
Rh001_022_018-    i_022    tia_h_in_001_018-    14854.152408945281
Rh001_023_018+    i_023    tia_h_in_001_018+    14828.43249241373
Rh001_023_018-    i_023    tia_h_in_001_018-    14549.153178843078
Rh001_024_018+    i_024    tia_h_in_001_018+    14697.54847242801
Rh001_024_018-    i_024    tia_h_in_001_018-    14738.329732505079
Rh001_025_018+    i_025    tia_h_in_001_018+    13938.575981854881
Rh001_025_018-    i_025    tia_h_in_001_018-    14931.930061381063
Rh001_026_018+    i_026    tia_h_in_001_018+    13084.866014029138
Rh001_026_018-    i_026    tia_h_in_001_018-    14965.12397122963
Rh001_027_018+    i_027    tia_h_in_001_018+    5000
Rh001_027_018-    i_027    tia_h_in_001_018-    14972.644783747533
Rh001_028_018+    i_028    tia_h_in_001_018+    13495.511678359035
Rh001_028_018-    i_028    tia_h_in_001_018-    15025.083306607119
Rh001_029_018+    i_029    tia_h_in_001_018+    14970.406232136895
Rh001_029_018-    i_029    tia_h_in_001_018-    13251.85473540874
Rh001_030_018+    i_030    tia_h_in_001_018+    15022.129646856009
Rh001_030_018-    i_030    tia_h_in_001_018-    12946.384727380064
Rh001_031_018+    i_031    tia_h_in_001_018+    13078.166114333
Rh001_031_018-    i_031    tia_h_in_001_018-    14957.444373791739
Rh001_032_018+    i_032    tia_h_in_001_018+    14964.770009514521
Rh001_032_018-    i_032    tia_h_in_001_018-    14734.006199598616
Rh001_033_018+    i_033    tia_h_in_001_018+    12335.057266905053
Rh001_033_018-    i_033    tia_h_in_001_018-    14869.740327654601
Rh001_034_018+    i_034    tia_h_in_001_018+    13592.486533191935
Rh001_034_018-    i_034    tia_h_in_001_018-    15123.86203365334
Rh001_035_018+    i_035    tia_h_in_001_018+    14951.814719904514
Rh001_035_018-    i_035    tia_h_in_001_018-    14364.761014990037
Rh001_036_018+    i_036    tia_h_in_001_018+    13928.696565152435
Rh001_036_018-    i_036    tia_h_in_001_018-    15128.727382248133
Rh001_037_018+    i_037    tia_h_in_001_018+    15000
Rh001_037_018-    i_037    tia_h_in_001_018-    15100.599208347825
Rh001_038_018+    i_038    tia_h_in_001_018+    13280.432276414072
Rh001_038_018-    i_038    tia_h_in_001_018-    15000
Rh001_039_018+    i_039    tia_h_in_001_018+    14068.888669262953
Rh001_039_018-    i_039    tia_h_in_001_018-    15081.389367701257
Rh001_040_018+    i_040    tia_h_in_001_018+    10882.577684548703
Rh001_040_018-    i_040    tia_h_in_001_018-    14823.27051352108
Rh001_041_018+    i_041    tia_h_in_001_018+    14922.38118989105
Rh001_041_018-    i_041    tia_h_in_001_018-    14369.940851465059
Rh001_042_018+    i_042    tia_h_in_001_018+    14956.184056943162
Rh001_042_018-    i_042    tia_h_in_001_018-    13814.998178536796
Rh001_043_018+    i_043    tia_h_in_001_018+    14943.018860150049
Rh001_043_018-    i_043    tia_h_in_001_018-    14621.80420021986
Rh001_044_018+    i_044    tia_h_in_001_018+    14791.797232462954
Rh001_044_018-    i_044    tia_h_in_001_018-    15036.378378609339
Rh001_045_018+    i_045    tia_h_in_001_018+    14892.395258592793
Rh001_045_018-    i_045    tia_h_in_001_018-    14514.54384478745
Rh001_046_018+    i_046    tia_h_in_001_018+    12211.331254490287
Rh001_046_018-    i_046    tia_h_in_001_018-    5000
Rh001_047_018+    i_047    tia_h_in_001_018+    13115.814906363574
Rh001_047_018-    i_047    tia_h_in_001_018-    15030.587545512628
Rh001_048_018+    i_048    tia_h_in_001_018+    12348.792021273932
Rh001_048_018-    i_048    tia_h_in_001_018-    14952.92237283507
Rh001_049_018+    i_049    tia_h_in_001_018+    14799.482761476182
Rh001_049_018-    i_049    tia_h_in_001_018-    14597.68153651466
Rh001_050_018+    i_050    tia_h_in_001_018+    14775.408643763869
Rh001_050_018-    i_050    tia_h_in_001_018-    15117.638966187493
Rh001_051_018+    i_051    tia_h_in_001_018+    14927.504152014375
Rh001_051_018-    i_051    tia_h_in_001_018-    14580.350238922156
Rh001_052_018+    i_052    tia_h_in_001_018+    15027.086350304879
Rh001_052_018-    i_052    tia_h_in_001_018-    14119.88740560564
Rh001_053_018+    i_053    tia_h_in_001_018+    15070.021978772213
Rh001_053_018-    i_053    tia_h_in_001_018-    14435.73328561633
Rh001_054_018+    i_054    tia_h_in_001_018+    14826.25875669571
Rh001_054_018-    i_054    tia_h_in_001_018-    13908.603177197887
Rh001_055_018+    i_055    tia_h_in_001_018+    14176.722496184559
Rh001_055_018-    i_055    tia_h_in_001_018-    14832.802727341827
Rh001_056_018+    i_056    tia_h_in_001_018+    15201.83728417483
Rh001_056_018-    i_056    tia_h_in_001_018-    10769.964998021334
Rh001_057_018+    i_057    tia_h_in_001_018+    13939.278223384947
Rh001_057_018-    i_057    tia_h_in_001_018-    5000
Rh001_058_018+    i_058    tia_h_in_001_018+    14646.264450778508
Rh001_058_018-    i_058    tia_h_in_001_018-    15174.889169806924
Rh001_059_018+    i_059    tia_h_in_001_018+    14879.54123784515
Rh001_059_018-    i_059    tia_h_in_001_018-    14331.941686156464
Rh001_060_018+    i_060    tia_h_in_001_018+    13005.674699664225
Rh001_060_018-    i_060    tia_h_in_001_018-    14795.774688293703
Rh001_061_018+    i_061    tia_h_in_001_018+    15093.26930612034
Rh001_061_018-    i_061    tia_h_in_001_018-    14200.1493942918
Rh001_062_018+    i_062    tia_h_in_001_018+    15081.637422574806
Rh001_062_018-    i_062    tia_h_in_001_018-    13326.443093312497
Rh001_063_018+    i_063    tia_h_in_001_018+    15161.73341412497
Rh001_063_018-    i_063    tia_h_in_001_018-    9874.442810918792
Rh001_064_018+    i_064    tia_h_in_001_018+    5000
Rh001_064_018-    i_064    tia_h_in_001_018-    11036.352166229004

* Neuron 19
Rh001_001_019+    i_001    tia_h_in_001_019+    15000
Rh001_001_019-    i_001    tia_h_in_001_019-    15103.970279272731
Rh001_002_019+    i_002    tia_h_in_001_019+    13323.852672635365
Rh001_002_019-    i_002    tia_h_in_001_019-    14935.321691588833
Rh001_003_019+    i_003    tia_h_in_001_019+    10621.699435462813
Rh001_003_019-    i_003    tia_h_in_001_019-    15075.465029655528
Rh001_004_019+    i_004    tia_h_in_001_019+    14289.647139229979
Rh001_004_019-    i_004    tia_h_in_001_019-    15148.048098833873
Rh001_005_019+    i_005    tia_h_in_001_019+    15129.519768511642
Rh001_005_019-    i_005    tia_h_in_001_019-    12824.750293537829
Rh001_006_019+    i_006    tia_h_in_001_019+    15000
Rh001_006_019-    i_006    tia_h_in_001_019-    11875.08010498886
Rh001_007_019+    i_007    tia_h_in_001_019+    15000
Rh001_007_019-    i_007    tia_h_in_001_019-    15000
Rh001_008_019+    i_008    tia_h_in_001_019+    14798.08254559627
Rh001_008_019-    i_008    tia_h_in_001_019-    12842.270179269934
Rh001_009_019+    i_009    tia_h_in_001_019+    14174.81625064668
Rh001_009_019-    i_009    tia_h_in_001_019-    15025.902004975562
Rh001_010_019+    i_010    tia_h_in_001_019+    12713.995513747379
Rh001_010_019-    i_010    tia_h_in_001_019-    15001.555590236656
Rh001_011_019+    i_011    tia_h_in_001_019+    14925.488111455288
Rh001_011_019-    i_011    tia_h_in_001_019-    14094.514815024635
Rh001_012_019+    i_012    tia_h_in_001_019+    14951.448673963205
Rh001_012_019-    i_012    tia_h_in_001_019-    5000
Rh001_013_019+    i_013    tia_h_in_001_019+    14972.348795128792
Rh001_013_019-    i_013    tia_h_in_001_019-    13252.744044858267
Rh001_014_019+    i_014    tia_h_in_001_019+    14924.522135033396
Rh001_014_019-    i_014    tia_h_in_001_019-    14362.868831096042
Rh001_015_019+    i_015    tia_h_in_001_019+    15044.958769474231
Rh001_015_019-    i_015    tia_h_in_001_019-    13991.770059868888
Rh001_016_019+    i_016    tia_h_in_001_019+    14141.129575849798
Rh001_016_019-    i_016    tia_h_in_001_019-    14912.860431164245
Rh001_017_019+    i_017    tia_h_in_001_019+    12158.527555733926
Rh001_017_019-    i_017    tia_h_in_001_019-    15000
Rh001_018_019+    i_018    tia_h_in_001_019+    12226.439141807065
Rh001_018_019-    i_018    tia_h_in_001_019-    14810.156221462446
Rh001_019_019+    i_019    tia_h_in_001_019+    14376.919383092214
Rh001_019_019-    i_019    tia_h_in_001_019-    14941.109232642757
Rh001_020_019+    i_020    tia_h_in_001_019+    14820.2017155839
Rh001_020_019-    i_020    tia_h_in_001_019-    14805.813208709314
Rh001_021_019+    i_021    tia_h_in_001_019+    14840.073543005909
Rh001_021_019-    i_021    tia_h_in_001_019-    13682.934415153763
Rh001_022_019+    i_022    tia_h_in_001_019+    15133.22633005557
Rh001_022_019-    i_022    tia_h_in_001_019-    14046.505250985696
Rh001_023_019+    i_023    tia_h_in_001_019+    14725.131907304869
Rh001_023_019-    i_023    tia_h_in_001_019-    15098.274542402745
Rh001_024_019+    i_024    tia_h_in_001_019+    14168.928798905108
Rh001_024_019-    i_024    tia_h_in_001_019-    14875.221168669766
Rh001_025_019+    i_025    tia_h_in_001_019+    12594.821637648762
Rh001_025_019-    i_025    tia_h_in_001_019-    15084.873588179309
Rh001_026_019+    i_026    tia_h_in_001_019+    5000
Rh001_026_019-    i_026    tia_h_in_001_019-    5000
Rh001_027_019+    i_027    tia_h_in_001_019+    14897.065807452325
Rh001_027_019-    i_027    tia_h_in_001_019-    13461.074920883788
Rh001_028_019+    i_028    tia_h_in_001_019+    15100.560512089594
Rh001_028_019-    i_028    tia_h_in_001_019-    14486.157870282792
Rh001_029_019+    i_029    tia_h_in_001_019+    15168.171786248393
Rh001_029_019-    i_029    tia_h_in_001_019-    13469.146529580683
Rh001_030_019+    i_030    tia_h_in_001_019+    15103.98353363744
Rh001_030_019-    i_030    tia_h_in_001_019-    13404.726332907661
Rh001_031_019+    i_031    tia_h_in_001_019+    13930.751293223428
Rh001_031_019-    i_031    tia_h_in_001_019-    15223.87493510029
Rh001_032_019+    i_032    tia_h_in_001_019+    13569.095924550653
Rh001_032_019-    i_032    tia_h_in_001_019-    14932.032408579433
Rh001_033_019+    i_033    tia_h_in_001_019+    13962.956004126525
Rh001_033_019-    i_033    tia_h_in_001_019-    15080.692450614857
Rh001_034_019+    i_034    tia_h_in_001_019+    14341.871816620542
Rh001_034_019-    i_034    tia_h_in_001_019-    15197.646320184187
Rh001_035_019+    i_035    tia_h_in_001_019+    14830.513526872788
Rh001_035_019-    i_035    tia_h_in_001_019-    13855.30147693797
Rh001_036_019+    i_036    tia_h_in_001_019+    15106.54447225725
Rh001_036_019-    i_036    tia_h_in_001_019-    13366.868402734735
Rh001_037_019+    i_037    tia_h_in_001_019+    5000
Rh001_037_019-    i_037    tia_h_in_001_019-    13245.280600952143
Rh001_038_019+    i_038    tia_h_in_001_019+    13856.013482238679
Rh001_038_019-    i_038    tia_h_in_001_019-    14942.574312511311
Rh001_039_019+    i_039    tia_h_in_001_019+    15120.559764992044
Rh001_039_019-    i_039    tia_h_in_001_019-    14866.142580486941
Rh001_040_019+    i_040    tia_h_in_001_019+    13128.016595191191
Rh001_040_019-    i_040    tia_h_in_001_019-    15012.631333355124
Rh001_041_019+    i_041    tia_h_in_001_019+    15112.996458334048
Rh001_041_019-    i_041    tia_h_in_001_019-    13506.467761893322
Rh001_042_019+    i_042    tia_h_in_001_019+    15046.276911544386
Rh001_042_019-    i_042    tia_h_in_001_019-    15000
Rh001_043_019+    i_043    tia_h_in_001_019+    15260.990303767421
Rh001_043_019-    i_043    tia_h_in_001_019-    12934.624489610227
Rh001_044_019+    i_044    tia_h_in_001_019+    14952.692384788263
Rh001_044_019-    i_044    tia_h_in_001_019-    14926.272587073461
Rh001_045_019+    i_045    tia_h_in_001_019+    5000
Rh001_045_019-    i_045    tia_h_in_001_019-    15049.171799974285
Rh001_046_019+    i_046    tia_h_in_001_019+    12533.003115323716
Rh001_046_019-    i_046    tia_h_in_001_019-    15020.505812705596
Rh001_047_019+    i_047    tia_h_in_001_019+    14044.46724831657
Rh001_047_019-    i_047    tia_h_in_001_019-    14978.415900024624
Rh001_048_019+    i_048    tia_h_in_001_019+    14046.717962742418
Rh001_048_019-    i_048    tia_h_in_001_019-    14975.730442434846
Rh001_049_019+    i_049    tia_h_in_001_019+    14961.741661788501
Rh001_049_019-    i_049    tia_h_in_001_019-    13360.780708451819
Rh001_050_019+    i_050    tia_h_in_001_019+    14773.013026548242
Rh001_050_019-    i_050    tia_h_in_001_019-    12970.549851548001
Rh001_051_019+    i_051    tia_h_in_001_019+    14912.098260509147
Rh001_051_019-    i_051    tia_h_in_001_019-    13058.114252838823
Rh001_052_019+    i_052    tia_h_in_001_019+    14853.661468233046
Rh001_052_019-    i_052    tia_h_in_001_019-    14878.68601800549
Rh001_053_019+    i_053    tia_h_in_001_019+    14989.251815674897
Rh001_053_019-    i_053    tia_h_in_001_019-    14822.642362092902
Rh001_054_019+    i_054    tia_h_in_001_019+    13001.577502032686
Rh001_054_019-    i_054    tia_h_in_001_019-    14938.421899231982
Rh001_055_019+    i_055    tia_h_in_001_019+    12137.11699974609
Rh001_055_019-    i_055    tia_h_in_001_019-    14971.249725469363
Rh001_056_019+    i_056    tia_h_in_001_019+    15047.05489945265
Rh001_056_019-    i_056    tia_h_in_001_019-    14916.638050016827
Rh001_057_019+    i_057    tia_h_in_001_019+    15105.78731479467
Rh001_057_019-    i_057    tia_h_in_001_019-    10683.17136683689
Rh001_058_019+    i_058    tia_h_in_001_019+    14868.746023313082
Rh001_058_019-    i_058    tia_h_in_001_019-    12914.810683943499
Rh001_059_019+    i_059    tia_h_in_001_019+    14841.379461173772
Rh001_059_019-    i_059    tia_h_in_001_019-    14350.304095999936
Rh001_060_019+    i_060    tia_h_in_001_019+    11432.607797243978
Rh001_060_019-    i_060    tia_h_in_001_019-    15264.629983587503
Rh001_061_019+    i_061    tia_h_in_001_019+    9842.651198769201
Rh001_061_019-    i_061    tia_h_in_001_019-    14800.078742797137
Rh001_062_019+    i_062    tia_h_in_001_019+    11756.474542063508
Rh001_062_019-    i_062    tia_h_in_001_019-    14893.431719681346
Rh001_063_019+    i_063    tia_h_in_001_019+    14857.329203008318
Rh001_063_019-    i_063    tia_h_in_001_019-    13548.380987736964
Rh001_064_019+    i_064    tia_h_in_001_019+    14901.42286750279
Rh001_064_019-    i_064    tia_h_in_001_019-    15000

* Neuron 20
Rh001_001_020+    i_001    tia_h_in_001_020+    14924.863017457405
Rh001_001_020-    i_001    tia_h_in_001_020-    13219.80965621961
Rh001_002_020+    i_002    tia_h_in_001_020+    15054.520886606833
Rh001_002_020-    i_002    tia_h_in_001_020-    12721.897712524322
Rh001_003_020+    i_003    tia_h_in_001_020+    15077.257322891053
Rh001_003_020-    i_003    tia_h_in_001_020-    12187.03295011494
Rh001_004_020+    i_004    tia_h_in_001_020+    5000
Rh001_004_020-    i_004    tia_h_in_001_020-    15045.811685102159
Rh001_005_020+    i_005    tia_h_in_001_020+    14949.737536169461
Rh001_005_020-    i_005    tia_h_in_001_020-    5000
Rh001_006_020+    i_006    tia_h_in_001_020+    13815.004870505421
Rh001_006_020-    i_006    tia_h_in_001_020-    15000
Rh001_007_020+    i_007    tia_h_in_001_020+    12934.128792308647
Rh001_007_020-    i_007    tia_h_in_001_020-    14906.057063780572
Rh001_008_020+    i_008    tia_h_in_001_020+    12919.421658023748
Rh001_008_020-    i_008    tia_h_in_001_020-    14980.474098978788
Rh001_009_020+    i_009    tia_h_in_001_020+    14812.887142798927
Rh001_009_020-    i_009    tia_h_in_001_020-    14772.780233003125
Rh001_010_020+    i_010    tia_h_in_001_020+    14931.358821129648
Rh001_010_020-    i_010    tia_h_in_001_020-    11383.77747704574
Rh001_011_020+    i_011    tia_h_in_001_020+    12091.634415388604
Rh001_011_020-    i_011    tia_h_in_001_020-    15000
Rh001_012_020+    i_012    tia_h_in_001_020+    12559.559444943545
Rh001_012_020-    i_012    tia_h_in_001_020-    15074.47814890298
Rh001_013_020+    i_013    tia_h_in_001_020+    15320.926397430092
Rh001_013_020-    i_013    tia_h_in_001_020-    14565.660027864742
Rh001_014_020+    i_014    tia_h_in_001_020+    12816.64328906838
Rh001_014_020-    i_014    tia_h_in_001_020-    15116.69486090714
Rh001_015_020+    i_015    tia_h_in_001_020+    14465.125587017534
Rh001_015_020-    i_015    tia_h_in_001_020-    14902.086550071379
Rh001_016_020+    i_016    tia_h_in_001_020+    5000
Rh001_016_020-    i_016    tia_h_in_001_020-    15172.599943841631
Rh001_017_020+    i_017    tia_h_in_001_020+    15067.93243333709
Rh001_017_020-    i_017    tia_h_in_001_020-    12120.51900037419
Rh001_018_020+    i_018    tia_h_in_001_020+    14169.86376353684
Rh001_018_020-    i_018    tia_h_in_001_020-    14700.74790954248
Rh001_019_020+    i_019    tia_h_in_001_020+    13808.909030720042
Rh001_019_020-    i_019    tia_h_in_001_020-    15144.266686041414
Rh001_020_020+    i_020    tia_h_in_001_020+    13650.08300098515
Rh001_020_020-    i_020    tia_h_in_001_020-    15021.726772884937
Rh001_021_020+    i_021    tia_h_in_001_020+    14930.980554349822
Rh001_021_020-    i_021    tia_h_in_001_020-    14487.267664227862
Rh001_022_020+    i_022    tia_h_in_001_020+    15166.7238131211
Rh001_022_020-    i_022    tia_h_in_001_020-    14218.12666421145
Rh001_023_020+    i_023    tia_h_in_001_020+    14710.592084748023
Rh001_023_020-    i_023    tia_h_in_001_020-    15219.578520564124
Rh001_024_020+    i_024    tia_h_in_001_020+    13072.808044646128
Rh001_024_020-    i_024    tia_h_in_001_020-    15056.401111913186
Rh001_025_020+    i_025    tia_h_in_001_020+    14801.400263000196
Rh001_025_020-    i_025    tia_h_in_001_020-    5000
Rh001_026_020+    i_026    tia_h_in_001_020+    14913.163634519266
Rh001_026_020-    i_026    tia_h_in_001_020-    15115.001410339348
Rh001_027_020+    i_027    tia_h_in_001_020+    14996.549598728367
Rh001_027_020-    i_027    tia_h_in_001_020-    14363.298405017085
Rh001_028_020+    i_028    tia_h_in_001_020+    15043.018891179932
Rh001_028_020-    i_028    tia_h_in_001_020-    12493.931365989372
Rh001_029_020+    i_029    tia_h_in_001_020+    14821.95706231133
Rh001_029_020-    i_029    tia_h_in_001_020-    13707.771009476768
Rh001_030_020+    i_030    tia_h_in_001_020+    14949.352010051394
Rh001_030_020-    i_030    tia_h_in_001_020-    14181.897407068624
Rh001_031_020+    i_031    tia_h_in_001_020+    14963.696133794703
Rh001_031_020-    i_031    tia_h_in_001_020-    13833.798224489736
Rh001_032_020+    i_032    tia_h_in_001_020+    14830.145465949143
Rh001_032_020-    i_032    tia_h_in_001_020-    15051.155656246472
Rh001_033_020+    i_033    tia_h_in_001_020+    14846.567725259181
Rh001_033_020-    i_033    tia_h_in_001_020-    15095.551739129745
Rh001_034_020+    i_034    tia_h_in_001_020+    15221.61254745699
Rh001_034_020-    i_034    tia_h_in_001_020-    14490.68604928724
Rh001_035_020+    i_035    tia_h_in_001_020+    15000
Rh001_035_020-    i_035    tia_h_in_001_020-    14892.492782755311
Rh001_036_020+    i_036    tia_h_in_001_020+    15030.734073217294
Rh001_036_020-    i_036    tia_h_in_001_020-    13816.419932772382
Rh001_037_020+    i_037    tia_h_in_001_020+    14954.08053110027
Rh001_037_020-    i_037    tia_h_in_001_020-    13281.507050465101
Rh001_038_020+    i_038    tia_h_in_001_020+    14312.31536403001
Rh001_038_020-    i_038    tia_h_in_001_020-    15141.626848825832
Rh001_039_020+    i_039    tia_h_in_001_020+    14175.743934463753
Rh001_039_020-    i_039    tia_h_in_001_020-    14877.341909401444
Rh001_040_020+    i_040    tia_h_in_001_020+    15227.075127480544
Rh001_040_020-    i_040    tia_h_in_001_020-    13437.923902242539
Rh001_041_020+    i_041    tia_h_in_001_020+    14693.774195331122
Rh001_041_020-    i_041    tia_h_in_001_020-    5000
Rh001_042_020+    i_042    tia_h_in_001_020+    5000
Rh001_042_020-    i_042    tia_h_in_001_020-    14951.770469050247
Rh001_043_020+    i_043    tia_h_in_001_020+    15013.372264338284
Rh001_043_020-    i_043    tia_h_in_001_020-    12471.067755923208
Rh001_044_020+    i_044    tia_h_in_001_020+    14967.987850097938
Rh001_044_020-    i_044    tia_h_in_001_020-    13146.878944160193
Rh001_045_020+    i_045    tia_h_in_001_020+    15000
Rh001_045_020-    i_045    tia_h_in_001_020-    15144.050549367517
Rh001_046_020+    i_046    tia_h_in_001_020+    13308.621699022928
Rh001_046_020-    i_046    tia_h_in_001_020-    15173.027312450307
Rh001_047_020+    i_047    tia_h_in_001_020+    13556.62569159711
Rh001_047_020-    i_047    tia_h_in_001_020-    14868.016375601163
Rh001_048_020+    i_048    tia_h_in_001_020+    14815.175327443221
Rh001_048_020-    i_048    tia_h_in_001_020-    14776.809783594888
Rh001_049_020+    i_049    tia_h_in_001_020+    13516.28581456472
Rh001_049_020-    i_049    tia_h_in_001_020-    5000
Rh001_050_020+    i_050    tia_h_in_001_020+    5000
Rh001_050_020-    i_050    tia_h_in_001_020-    14858.810955676447
Rh001_051_020+    i_051    tia_h_in_001_020+    12875.426211547143
Rh001_051_020-    i_051    tia_h_in_001_020-    15080.364243849293
Rh001_052_020+    i_052    tia_h_in_001_020+    13647.174249654641
Rh001_052_020-    i_052    tia_h_in_001_020-    14970.603502814522
Rh001_053_020+    i_053    tia_h_in_001_020+    14499.059831472132
Rh001_053_020-    i_053    tia_h_in_001_020-    15000
Rh001_054_020+    i_054    tia_h_in_001_020+    13556.418290136138
Rh001_054_020-    i_054    tia_h_in_001_020-    15003.995277023196
Rh001_055_020+    i_055    tia_h_in_001_020+    14992.975705231034
Rh001_055_020-    i_055    tia_h_in_001_020-    12078.663439006637
Rh001_056_020+    i_056    tia_h_in_001_020+    15150.286568831256
Rh001_056_020-    i_056    tia_h_in_001_020-    14351.369827188733
Rh001_057_020+    i_057    tia_h_in_001_020+    13231.916501133102
Rh001_057_020-    i_057    tia_h_in_001_020-    15000
Rh001_058_020+    i_058    tia_h_in_001_020+    13891.63194689789
Rh001_058_020-    i_058    tia_h_in_001_020-    15040.143121527677
Rh001_059_020+    i_059    tia_h_in_001_020+    12584.09664318536
Rh001_059_020-    i_059    tia_h_in_001_020-    15208.023528248073
Rh001_060_020+    i_060    tia_h_in_001_020+    14670.387656700968
Rh001_060_020-    i_060    tia_h_in_001_020-    15076.631175825616
Rh001_061_020+    i_061    tia_h_in_001_020+    14797.770681696364
Rh001_061_020-    i_061    tia_h_in_001_020-    15000
Rh001_062_020+    i_062    tia_h_in_001_020+    14980.871963286218
Rh001_062_020-    i_062    tia_h_in_001_020-    12297.433177920373
Rh001_063_020+    i_063    tia_h_in_001_020+    14982.961901137209
Rh001_063_020-    i_063    tia_h_in_001_020-    11509.976092666839
Rh001_064_020+    i_064    tia_h_in_001_020+    15034.804018878567
Rh001_064_020-    i_064    tia_h_in_001_020-    15000

* ----- Bias
    
        
Rb_h001_001+    b_001    tia_h_in_001_001+    15078.395532925888
Rb_h001_001-    b_001    tia_h_in_001_001-    15000
Rb_h001_002+    b_001    tia_h_in_001_002+    11872.443048221114
Rb_h001_002-    b_001    tia_h_in_001_002-    15054.46664406758
Rb_h001_003+    b_001    tia_h_in_001_003+    15045.88856393484
Rb_h001_003-    b_001    tia_h_in_001_003-    9616.338244369168
Rb_h001_004+    b_001    tia_h_in_001_004+    15061.105093063703
Rb_h001_004-    b_001    tia_h_in_001_004-    13623.293416486838
Rb_h001_005+    b_001    tia_h_in_001_005+    5000
Rb_h001_005-    b_001    tia_h_in_001_005-    15079.764394366393
Rb_h001_006+    b_001    tia_h_in_001_006+    14377.910198733247
Rb_h001_006-    b_001    tia_h_in_001_006-    14918.846117493054
Rb_h001_007+    b_001    tia_h_in_001_007+    13200.892193227548
Rb_h001_007-    b_001    tia_h_in_001_007-    15093.480176814763
Rb_h001_008+    b_001    tia_h_in_001_008+    12912.975010181182
Rb_h001_008-    b_001    tia_h_in_001_008-    14896.008342822312
Rb_h001_009+    b_001    tia_h_in_001_009+    12150.995342167178
Rb_h001_009-    b_001    tia_h_in_001_009-    15162.95080775998
Rb_h001_010+    b_001    tia_h_in_001_010+    15110.272170555823
Rb_h001_010-    b_001    tia_h_in_001_010-    14305.114474490654
Rb_h001_011+    b_001    tia_h_in_001_011+    12290.018053493484
Rb_h001_011-    b_001    tia_h_in_001_011-    15022.78171971052
Rb_h001_012+    b_001    tia_h_in_001_012+    11437.596762624746
Rb_h001_012-    b_001    tia_h_in_001_012-    15042.024009009217
Rb_h001_013+    b_001    tia_h_in_001_013+    13821.211157765314
Rb_h001_013-    b_001    tia_h_in_001_013-    15075.945732327798
Rb_h001_014+    b_001    tia_h_in_001_014+    15108.713771909508
Rb_h001_014-    b_001    tia_h_in_001_014-    13705.821830965895
Rb_h001_015+    b_001    tia_h_in_001_015+    15000
Rb_h001_015-    b_001    tia_h_in_001_015-    15070.496020153065
Rb_h001_016+    b_001    tia_h_in_001_016+    15013.386519462485
Rb_h001_016-    b_001    tia_h_in_001_016-    12250.421471499283
Rb_h001_017+    b_001    tia_h_in_001_017+    15092.315641328198
Rb_h001_017-    b_001    tia_h_in_001_017-    13123.843828451403
Rb_h001_018+    b_001    tia_h_in_001_018+    5000
Rb_h001_018-    b_001    tia_h_in_001_018-    15140.532525137914
Rb_h001_019+    b_001    tia_h_in_001_019+    14937.270178482904
Rb_h001_019-    b_001    tia_h_in_001_019-    9532.130610346165
Rb_h001_020+    b_001    tia_h_in_001_020+    11799.25518286704
Rb_h001_020-    b_001    tia_h_in_001_020-    15175.697662556679

* ----- Weights
* Layer 002

* Neuron 1
Rh002_001_001+    hidden_activ_out_h001_001    tia_h_in_002_001+    5000
Rh002_001_001-    hidden_activ_out_h001_001    tia_h_in_002_001-    6456.253518247686
Rh002_002_001+    hidden_activ_out_h001_002    tia_h_in_002_001+    5000
Rh002_002_001-    hidden_activ_out_h001_002    tia_h_in_002_001-    15037.151548310534
Rh002_003_001+    hidden_activ_out_h001_003    tia_h_in_002_001+    14881.471927053644
Rh002_003_001-    hidden_activ_out_h001_003    tia_h_in_002_001-    6422.7945025988065
Rh002_004_001+    hidden_activ_out_h001_004    tia_h_in_002_001+    5000
Rh002_004_001-    hidden_activ_out_h001_004    tia_h_in_002_001-    13096.608028316716
Rh002_005_001+    hidden_activ_out_h001_005    tia_h_in_002_001+    5712.847520661422
Rh002_005_001-    hidden_activ_out_h001_005    tia_h_in_002_001-    15210.213140433552
Rh002_006_001+    hidden_activ_out_h001_006    tia_h_in_002_001+    15098.051709243735
Rh002_006_001-    hidden_activ_out_h001_006    tia_h_in_002_001-    14941.978189431404
Rh002_007_001+    hidden_activ_out_h001_007    tia_h_in_002_001+    11576.471285291558
Rh002_007_001-    hidden_activ_out_h001_007    tia_h_in_002_001-    14986.203209317562
Rh002_008_001+    hidden_activ_out_h001_008    tia_h_in_002_001+    5946.043018467675
Rh002_008_001-    hidden_activ_out_h001_008    tia_h_in_002_001-    15140.377491096613
Rh002_009_001+    hidden_activ_out_h001_009    tia_h_in_002_001+    10412.552503349454
Rh002_009_001-    hidden_activ_out_h001_009    tia_h_in_002_001-    14955.63894360923
Rh002_010_001+    hidden_activ_out_h001_010    tia_h_in_002_001+    15174.58299863723
Rh002_010_001-    hidden_activ_out_h001_010    tia_h_in_002_001-    14403.143306301883
Rh002_011_001+    hidden_activ_out_h001_011    tia_h_in_002_001+    8286.202376542484
Rh002_011_001-    hidden_activ_out_h001_011    tia_h_in_002_001-    14886.090605850568
Rh002_012_001+    hidden_activ_out_h001_012    tia_h_in_002_001+    15111.579409798329
Rh002_012_001-    hidden_activ_out_h001_012    tia_h_in_002_001-    5000
Rh002_013_001+    hidden_activ_out_h001_013    tia_h_in_002_001+    8366.634085386013
Rh002_013_001-    hidden_activ_out_h001_013    tia_h_in_002_001-    15086.206553509755
Rh002_014_001+    hidden_activ_out_h001_014    tia_h_in_002_001+    15364.257959553033
Rh002_014_001-    hidden_activ_out_h001_014    tia_h_in_002_001-    14935.72696662942
Rh002_015_001+    hidden_activ_out_h001_015    tia_h_in_002_001+    14965.7011496528
Rh002_015_001-    hidden_activ_out_h001_015    tia_h_in_002_001-    15000
Rh002_016_001+    hidden_activ_out_h001_016    tia_h_in_002_001+    15028.858155226984
Rh002_016_001-    hidden_activ_out_h001_016    tia_h_in_002_001-    7064.22445054274
Rh002_017_001+    hidden_activ_out_h001_017    tia_h_in_002_001+    15135.672465922624
Rh002_017_001-    hidden_activ_out_h001_017    tia_h_in_002_001-    6646.114434545529
Rh002_018_001+    hidden_activ_out_h001_018    tia_h_in_002_001+    11960.062432188039
Rh002_018_001-    hidden_activ_out_h001_018    tia_h_in_002_001-    14940.305928450543
Rh002_019_001+    hidden_activ_out_h001_019    tia_h_in_002_001+    15083.303482433757
Rh002_019_001-    hidden_activ_out_h001_019    tia_h_in_002_001-    6003.496666427148
Rh002_020_001+    hidden_activ_out_h001_020    tia_h_in_002_001+    15120.337432251146
Rh002_020_001-    hidden_activ_out_h001_020    tia_h_in_002_001-    15000

* Neuron 2
Rh002_001_002+    hidden_activ_out_h001_001    tia_h_in_002_002+    14999.60969178854
Rh002_001_002-    hidden_activ_out_h001_001    tia_h_in_002_002-    11825.413162083463
Rh002_002_002+    hidden_activ_out_h001_002    tia_h_in_002_002+    14986.803736677717
Rh002_002_002-    hidden_activ_out_h001_002    tia_h_in_002_002-    15000
Rh002_003_002+    hidden_activ_out_h001_003    tia_h_in_002_002+    10067.170492432635
Rh002_003_002-    hidden_activ_out_h001_003    tia_h_in_002_002-    15083.557637066791
Rh002_004_002+    hidden_activ_out_h001_004    tia_h_in_002_002+    12947.756778254863
Rh002_004_002-    hidden_activ_out_h001_004    tia_h_in_002_002-    15099.211123512545
Rh002_005_002+    hidden_activ_out_h001_005    tia_h_in_002_002+    15040.22766420946
Rh002_005_002-    hidden_activ_out_h001_005    tia_h_in_002_002-    7884.478758276538
Rh002_006_002+    hidden_activ_out_h001_006    tia_h_in_002_002+    14276.614736654165
Rh002_006_002-    hidden_activ_out_h001_006    tia_h_in_002_002-    14769.595446190893
Rh002_007_002+    hidden_activ_out_h001_007    tia_h_in_002_002+    15155.477593718775
Rh002_007_002-    hidden_activ_out_h001_007    tia_h_in_002_002-    7335.2101238370615
Rh002_008_002+    hidden_activ_out_h001_008    tia_h_in_002_002+    15140.767276380055
Rh002_008_002-    hidden_activ_out_h001_008    tia_h_in_002_002-    7390.530168926109
Rh002_009_002+    hidden_activ_out_h001_009    tia_h_in_002_002+    14948.769341404157
Rh002_009_002-    hidden_activ_out_h001_009    tia_h_in_002_002-    7394.270508016872
Rh002_010_002+    hidden_activ_out_h001_010    tia_h_in_002_002+    13147.118199748049
Rh002_010_002-    hidden_activ_out_h001_010    tia_h_in_002_002-    14681.393773515676
Rh002_011_002+    hidden_activ_out_h001_011    tia_h_in_002_002+    15293.81895212824
Rh002_011_002-    hidden_activ_out_h001_011    tia_h_in_002_002-    7152.534343327828
Rh002_012_002+    hidden_activ_out_h001_012    tia_h_in_002_002+    15112.443067853277
Rh002_012_002-    hidden_activ_out_h001_012    tia_h_in_002_002-    9774.162305732047
Rh002_013_002+    hidden_activ_out_h001_013    tia_h_in_002_002+    15026.508198123773
Rh002_013_002-    hidden_activ_out_h001_013    tia_h_in_002_002-    6709.514329020705
Rh002_014_002+    hidden_activ_out_h001_014    tia_h_in_002_002+    15025.449817298468
Rh002_014_002-    hidden_activ_out_h001_014    tia_h_in_002_002-    14475.013068882536
Rh002_015_002+    hidden_activ_out_h001_015    tia_h_in_002_002+    12631.769660750035
Rh002_015_002-    hidden_activ_out_h001_015    tia_h_in_002_002-    14907.288004558988
Rh002_016_002+    hidden_activ_out_h001_016    tia_h_in_002_002+    14937.252725987553
Rh002_016_002-    hidden_activ_out_h001_016    tia_h_in_002_002-    15000
Rh002_017_002+    hidden_activ_out_h001_017    tia_h_in_002_002+    14728.084672464529
Rh002_017_002-    hidden_activ_out_h001_017    tia_h_in_002_002-    15121.816266606766
Rh002_018_002+    hidden_activ_out_h001_018    tia_h_in_002_002+    15147.968859187326
Rh002_018_002-    hidden_activ_out_h001_018    tia_h_in_002_002-    6638.207955342782
Rh002_019_002+    hidden_activ_out_h001_019    tia_h_in_002_002+    9652.921597792654
Rh002_019_002-    hidden_activ_out_h001_019    tia_h_in_002_002-    14968.741764470735
Rh002_020_002+    hidden_activ_out_h001_020    tia_h_in_002_002+    14745.92769091595
Rh002_020_002-    hidden_activ_out_h001_020    tia_h_in_002_002-    7966.534286456128

* Neuron 3
Rh002_001_003+    hidden_activ_out_h001_001    tia_h_in_002_003+    10124.130534824746
Rh002_001_003-    hidden_activ_out_h001_001    tia_h_in_002_003-    15009.626717456604
Rh002_002_003+    hidden_activ_out_h001_002    tia_h_in_002_003+    15055.901863971065
Rh002_002_003-    hidden_activ_out_h001_002    tia_h_in_002_003-    6446.786425168265
Rh002_003_003+    hidden_activ_out_h001_003    tia_h_in_002_003+    12250.106483401452
Rh002_003_003-    hidden_activ_out_h001_003    tia_h_in_002_003-    14950.982958267177
Rh002_004_003+    hidden_activ_out_h001_004    tia_h_in_002_003+    13997.086485952435
Rh002_004_003-    hidden_activ_out_h001_004    tia_h_in_002_003-    15128.817399961483
Rh002_005_003+    hidden_activ_out_h001_005    tia_h_in_002_003+    14988.224622740396
Rh002_005_003-    hidden_activ_out_h001_005    tia_h_in_002_003-    8828.797669697895
Rh002_006_003+    hidden_activ_out_h001_006    tia_h_in_002_003+    15214.32644164981
Rh002_006_003-    hidden_activ_out_h001_006    tia_h_in_002_003-    14592.04796029643
Rh002_007_003+    hidden_activ_out_h001_007    tia_h_in_002_003+    15091.289929841825
Rh002_007_003-    hidden_activ_out_h001_007    tia_h_in_002_003-    9586.3961934459
Rh002_008_003+    hidden_activ_out_h001_008    tia_h_in_002_003+    15005.944565623371
Rh002_008_003-    hidden_activ_out_h001_008    tia_h_in_002_003-    10327.3046915803
Rh002_009_003+    hidden_activ_out_h001_009    tia_h_in_002_003+    15273.567609369416
Rh002_009_003-    hidden_activ_out_h001_009    tia_h_in_002_003-    7934.166187204371
Rh002_010_003+    hidden_activ_out_h001_010    tia_h_in_002_003+    15027.751941287559
Rh002_010_003-    hidden_activ_out_h001_010    tia_h_in_002_003-    5000
Rh002_011_003+    hidden_activ_out_h001_011    tia_h_in_002_003+    15156.689123811433
Rh002_011_003-    hidden_activ_out_h001_011    tia_h_in_002_003-    8278.631043958023
Rh002_012_003+    hidden_activ_out_h001_012    tia_h_in_002_003+    15000
Rh002_012_003-    hidden_activ_out_h001_012    tia_h_in_002_003-    10738.90477718949
Rh002_013_003+    hidden_activ_out_h001_013    tia_h_in_002_003+    14941.35265803551
Rh002_013_003-    hidden_activ_out_h001_013    tia_h_in_002_003-    7905.450505881258
Rh002_014_003+    hidden_activ_out_h001_014    tia_h_in_002_003+    13207.34651040314
Rh002_014_003-    hidden_activ_out_h001_014    tia_h_in_002_003-    14916.24662396026
Rh002_015_003+    hidden_activ_out_h001_015    tia_h_in_002_003+    14658.223957063872
Rh002_015_003-    hidden_activ_out_h001_015    tia_h_in_002_003-    15082.673548952996
Rh002_016_003+    hidden_activ_out_h001_016    tia_h_in_002_003+    10411.047413235065
Rh002_016_003-    hidden_activ_out_h001_016    tia_h_in_002_003-    14954.766725608275
Rh002_017_003+    hidden_activ_out_h001_017    tia_h_in_002_003+    15025.364770812097
Rh002_017_003-    hidden_activ_out_h001_017    tia_h_in_002_003-    10065.747739010185
Rh002_018_003+    hidden_activ_out_h001_018    tia_h_in_002_003+    14931.166379513605
Rh002_018_003-    hidden_activ_out_h001_018    tia_h_in_002_003-    9995.030642405165
Rh002_019_003+    hidden_activ_out_h001_019    tia_h_in_002_003+    13019.46955146768
Rh002_019_003-    hidden_activ_out_h001_019    tia_h_in_002_003-    15264.990396608016
Rh002_020_003+    hidden_activ_out_h001_020    tia_h_in_002_003+    14989.536629710467
Rh002_020_003-    hidden_activ_out_h001_020    tia_h_in_002_003-    12095.32255229942

* Neuron 4
Rh002_001_004+    hidden_activ_out_h001_001    tia_h_in_002_004+    15000
Rh002_001_004-    hidden_activ_out_h001_001    tia_h_in_002_004-    15088.004923492852
Rh002_002_004+    hidden_activ_out_h001_002    tia_h_in_002_004+    15012.019609195506
Rh002_002_004-    hidden_activ_out_h001_002    tia_h_in_002_004-    10476.507282658475
Rh002_003_004+    hidden_activ_out_h001_003    tia_h_in_002_004+    10929.96384895176
Rh002_003_004-    hidden_activ_out_h001_003    tia_h_in_002_004-    15017.053105755891
Rh002_004_004+    hidden_activ_out_h001_004    tia_h_in_002_004+    14963.177079003659
Rh002_004_004-    hidden_activ_out_h001_004    tia_h_in_002_004-    13054.442098020843
Rh002_005_004+    hidden_activ_out_h001_005    tia_h_in_002_004+    15042.060139754873
Rh002_005_004-    hidden_activ_out_h001_005    tia_h_in_002_004-    9659.986948559317
Rh002_006_004+    hidden_activ_out_h001_006    tia_h_in_002_004+    5000
Rh002_006_004-    hidden_activ_out_h001_006    tia_h_in_002_004-    14874.2077082753
Rh002_007_004+    hidden_activ_out_h001_007    tia_h_in_002_004+    14785.251679409677
Rh002_007_004-    hidden_activ_out_h001_007    tia_h_in_002_004-    11550.626105162417
Rh002_008_004+    hidden_activ_out_h001_008    tia_h_in_002_004+    15094.385627334701
Rh002_008_004-    hidden_activ_out_h001_008    tia_h_in_002_004-    15000
Rh002_009_004+    hidden_activ_out_h001_009    tia_h_in_002_004+    15273.617286521383
Rh002_009_004-    hidden_activ_out_h001_009    tia_h_in_002_004-    13697.333146073162
Rh002_010_004+    hidden_activ_out_h001_010    tia_h_in_002_004+    15055.707671751388
Rh002_010_004-    hidden_activ_out_h001_010    tia_h_in_002_004-    12712.129333369861
Rh002_011_004+    hidden_activ_out_h001_011    tia_h_in_002_004+    15202.873608674034
Rh002_011_004-    hidden_activ_out_h001_011    tia_h_in_002_004-    11476.899590411855
Rh002_012_004+    hidden_activ_out_h001_012    tia_h_in_002_004+    14926.630622301956
Rh002_012_004-    hidden_activ_out_h001_012    tia_h_in_002_004-    5000
Rh002_013_004+    hidden_activ_out_h001_013    tia_h_in_002_004+    15039.028594513702
Rh002_013_004-    hidden_activ_out_h001_013    tia_h_in_002_004-    12164.539327591141
Rh002_014_004+    hidden_activ_out_h001_014    tia_h_in_002_004+    15041.284338107962
Rh002_014_004-    hidden_activ_out_h001_014    tia_h_in_002_004-    14329.440419105233
Rh002_015_004+    hidden_activ_out_h001_015    tia_h_in_002_004+    13089.61949343286
Rh002_015_004-    hidden_activ_out_h001_015    tia_h_in_002_004-    15113.777496545388
Rh002_016_004+    hidden_activ_out_h001_016    tia_h_in_002_004+    8770.529312197275
Rh002_016_004-    hidden_activ_out_h001_016    tia_h_in_002_004-    15007.209281912345
Rh002_017_004+    hidden_activ_out_h001_017    tia_h_in_002_004+    5000
Rh002_017_004-    hidden_activ_out_h001_017    tia_h_in_002_004-    15045.447363166424
Rh002_018_004+    hidden_activ_out_h001_018    tia_h_in_002_004+    15000
Rh002_018_004-    hidden_activ_out_h001_018    tia_h_in_002_004-    14192.210403285271
Rh002_019_004+    hidden_activ_out_h001_019    tia_h_in_002_004+    9439.399181001067
Rh002_019_004-    hidden_activ_out_h001_019    tia_h_in_002_004-    14887.390434032373
Rh002_020_004+    hidden_activ_out_h001_020    tia_h_in_002_004+    14882.531726566865
Rh002_020_004-    hidden_activ_out_h001_020    tia_h_in_002_004-    14701.941341207268

* Neuron 5
Rh002_001_005+    hidden_activ_out_h001_001    tia_h_in_002_005+    9520.650848771933
Rh002_001_005-    hidden_activ_out_h001_001    tia_h_in_002_005-    14947.436868697321
Rh002_002_005+    hidden_activ_out_h001_002    tia_h_in_002_005+    14983.871818746977
Rh002_002_005-    hidden_activ_out_h001_002    tia_h_in_002_005-    10361.345066967173
Rh002_003_005+    hidden_activ_out_h001_003    tia_h_in_002_005+    11769.551547306475
Rh002_003_005-    hidden_activ_out_h001_003    tia_h_in_002_005-    14917.261676838854
Rh002_004_005+    hidden_activ_out_h001_004    tia_h_in_002_005+    14385.090143403133
Rh002_004_005-    hidden_activ_out_h001_004    tia_h_in_002_005-    15124.738009422279
Rh002_005_005+    hidden_activ_out_h001_005    tia_h_in_002_005+    14997.877166584925
Rh002_005_005-    hidden_activ_out_h001_005    tia_h_in_002_005-    15000
Rh002_006_005+    hidden_activ_out_h001_006    tia_h_in_002_005+    14831.244895466312
Rh002_006_005-    hidden_activ_out_h001_006    tia_h_in_002_005-    12569.157002327078
Rh002_007_005+    hidden_activ_out_h001_007    tia_h_in_002_005+    14942.779072504843
Rh002_007_005-    hidden_activ_out_h001_007    tia_h_in_002_005-    11363.49443938834
Rh002_008_005+    hidden_activ_out_h001_008    tia_h_in_002_005+    14899.46501427033
Rh002_008_005-    hidden_activ_out_h001_008    tia_h_in_002_005-    10417.829970316441
Rh002_009_005+    hidden_activ_out_h001_009    tia_h_in_002_005+    14856.763485986652
Rh002_009_005-    hidden_activ_out_h001_009    tia_h_in_002_005-    13016.006414767997
Rh002_010_005+    hidden_activ_out_h001_010    tia_h_in_002_005+    14952.685500586464
Rh002_010_005-    hidden_activ_out_h001_010    tia_h_in_002_005-    14147.631862662385
Rh002_011_005+    hidden_activ_out_h001_011    tia_h_in_002_005+    14941.496649730834
Rh002_011_005-    hidden_activ_out_h001_011    tia_h_in_002_005-    5000
Rh002_012_005+    hidden_activ_out_h001_012    tia_h_in_002_005+    15039.899908774547
Rh002_012_005-    hidden_activ_out_h001_012    tia_h_in_002_005-    14417.243334764986
Rh002_013_005+    hidden_activ_out_h001_013    tia_h_in_002_005+    14872.326433111766
Rh002_013_005-    hidden_activ_out_h001_013    tia_h_in_002_005-    11833.453444279403
Rh002_014_005+    hidden_activ_out_h001_014    tia_h_in_002_005+    14524.59403513215
Rh002_014_005-    hidden_activ_out_h001_014    tia_h_in_002_005-    15177.970967694391
Rh002_015_005+    hidden_activ_out_h001_015    tia_h_in_002_005+    15137.884644687356
Rh002_015_005-    hidden_activ_out_h001_015    tia_h_in_002_005-    13296.826770307951
Rh002_016_005+    hidden_activ_out_h001_016    tia_h_in_002_005+    9679.664480239104
Rh002_016_005-    hidden_activ_out_h001_016    tia_h_in_002_005-    15149.219501930633
Rh002_017_005+    hidden_activ_out_h001_017    tia_h_in_002_005+    11556.193086341662
Rh002_017_005-    hidden_activ_out_h001_017    tia_h_in_002_005-    14997.76289137627
Rh002_018_005+    hidden_activ_out_h001_018    tia_h_in_002_005+    14941.951536099206
Rh002_018_005-    hidden_activ_out_h001_018    tia_h_in_002_005-    14017.566577731934
Rh002_019_005+    hidden_activ_out_h001_019    tia_h_in_002_005+    15000
Rh002_019_005-    hidden_activ_out_h001_019    tia_h_in_002_005-    14722.475347174288
Rh002_020_005+    hidden_activ_out_h001_020    tia_h_in_002_005+    14479.614366789217
Rh002_020_005-    hidden_activ_out_h001_020    tia_h_in_002_005-    14987.134996279525

* Neuron 6
Rh002_001_006+    hidden_activ_out_h001_001    tia_h_in_002_006+    14975.871651003094
Rh002_001_006-    hidden_activ_out_h001_001    tia_h_in_002_006-    15000
Rh002_002_006+    hidden_activ_out_h001_002    tia_h_in_002_006+    13022.881731441741
Rh002_002_006-    hidden_activ_out_h001_002    tia_h_in_002_006-    15095.265034346194
Rh002_003_006+    hidden_activ_out_h001_003    tia_h_in_002_006+    15152.010891727165
Rh002_003_006-    hidden_activ_out_h001_003    tia_h_in_002_006-    5675.071229752269
Rh002_004_006+    hidden_activ_out_h001_004    tia_h_in_002_006+    14898.131138385796
Rh002_004_006-    hidden_activ_out_h001_004    tia_h_in_002_006-    14689.194591551519
Rh002_005_006+    hidden_activ_out_h001_005    tia_h_in_002_006+    6175.927883905496
Rh002_005_006-    hidden_activ_out_h001_005    tia_h_in_002_006-    15091.006572837796
Rh002_006_006+    hidden_activ_out_h001_006    tia_h_in_002_006+    14828.434907386787
Rh002_006_006-    hidden_activ_out_h001_006    tia_h_in_002_006-    15114.660383399287
Rh002_007_006+    hidden_activ_out_h001_007    tia_h_in_002_006+    11325.083573419428
Rh002_007_006-    hidden_activ_out_h001_007    tia_h_in_002_006-    15031.829328372125
Rh002_008_006+    hidden_activ_out_h001_008    tia_h_in_002_006+    6694.078222393759
Rh002_008_006-    hidden_activ_out_h001_008    tia_h_in_002_006-    14718.28928227012
Rh002_009_006+    hidden_activ_out_h001_009    tia_h_in_002_006+    11796.113629904776
Rh002_009_006-    hidden_activ_out_h001_009    tia_h_in_002_006-    15169.654336356423
Rh002_010_006+    hidden_activ_out_h001_010    tia_h_in_002_006+    14919.441565730813
Rh002_010_006-    hidden_activ_out_h001_010    tia_h_in_002_006-    13678.156470117525
Rh002_011_006+    hidden_activ_out_h001_011    tia_h_in_002_006+    9367.630841163587
Rh002_011_006-    hidden_activ_out_h001_011    tia_h_in_002_006-    14895.434426150348
Rh002_012_006+    hidden_activ_out_h001_012    tia_h_in_002_006+    14920.107346909524
Rh002_012_006-    hidden_activ_out_h001_012    tia_h_in_002_006-    14077.111915924093
Rh002_013_006+    hidden_activ_out_h001_013    tia_h_in_002_006+    9334.276301717786
Rh002_013_006-    hidden_activ_out_h001_013    tia_h_in_002_006-    15054.267036491236
Rh002_014_006+    hidden_activ_out_h001_014    tia_h_in_002_006+    14580.898185736492
Rh002_014_006-    hidden_activ_out_h001_014    tia_h_in_002_006-    14896.164678158077
Rh002_015_006+    hidden_activ_out_h001_015    tia_h_in_002_006+    15130.022466309007
Rh002_015_006-    hidden_activ_out_h001_015    tia_h_in_002_006-    14848.60453000481
Rh002_016_006+    hidden_activ_out_h001_016    tia_h_in_002_006+    14816.148130157846
Rh002_016_006-    hidden_activ_out_h001_016    tia_h_in_002_006-    15000
Rh002_017_006+    hidden_activ_out_h001_017    tia_h_in_002_006+    5000
Rh002_017_006-    hidden_activ_out_h001_017    tia_h_in_002_006-    8565.166228227885
Rh002_018_006+    hidden_activ_out_h001_018    tia_h_in_002_006+    10331.256266528988
Rh002_018_006-    hidden_activ_out_h001_018    tia_h_in_002_006-    14924.114461156847
Rh002_019_006+    hidden_activ_out_h001_019    tia_h_in_002_006+    15099.029660866849
Rh002_019_006-    hidden_activ_out_h001_019    tia_h_in_002_006-    5122.738691994314
Rh002_020_006+    hidden_activ_out_h001_020    tia_h_in_002_006+    15047.404529560787
Rh002_020_006-    hidden_activ_out_h001_020    tia_h_in_002_006-    15000

* Neuron 7
Rh002_001_007+    hidden_activ_out_h001_001    tia_h_in_002_007+    11661.490726473046
Rh002_001_007-    hidden_activ_out_h001_001    tia_h_in_002_007-    15120.032446675606
Rh002_002_007+    hidden_activ_out_h001_002    tia_h_in_002_007+    15052.635014801053
Rh002_002_007-    hidden_activ_out_h001_002    tia_h_in_002_007-    7521.597049237151
Rh002_003_007+    hidden_activ_out_h001_003    tia_h_in_002_007+    15000
Rh002_003_007-    hidden_activ_out_h001_003    tia_h_in_002_007-    15084.552844947262
Rh002_004_007+    hidden_activ_out_h001_004    tia_h_in_002_007+    14935.955691734274
Rh002_004_007-    hidden_activ_out_h001_004    tia_h_in_002_007-    5000
Rh002_005_007+    hidden_activ_out_h001_005    tia_h_in_002_007+    14862.230094160217
Rh002_005_007-    hidden_activ_out_h001_005    tia_h_in_002_007-    15000
Rh002_006_007+    hidden_activ_out_h001_006    tia_h_in_002_007+    15193.393496638499
Rh002_006_007-    hidden_activ_out_h001_006    tia_h_in_002_007-    13938.73349364498
Rh002_007_007+    hidden_activ_out_h001_007    tia_h_in_002_007+    15023.376331727168
Rh002_007_007-    hidden_activ_out_h001_007    tia_h_in_002_007-    9361.8367481746
Rh002_008_007+    hidden_activ_out_h001_008    tia_h_in_002_007+    14958.820726974946
Rh002_008_007-    hidden_activ_out_h001_008    tia_h_in_002_007-    10262.377309544874
Rh002_009_007+    hidden_activ_out_h001_009    tia_h_in_002_007+    14888.351891680506
Rh002_009_007-    hidden_activ_out_h001_009    tia_h_in_002_007-    9460.538567476007
Rh002_010_007+    hidden_activ_out_h001_010    tia_h_in_002_007+    12697.24856146023
Rh002_010_007-    hidden_activ_out_h001_010    tia_h_in_002_007-    15032.400585226242
Rh002_011_007+    hidden_activ_out_h001_011    tia_h_in_002_007+    15223.875876196567
Rh002_011_007-    hidden_activ_out_h001_011    tia_h_in_002_007-    8442.427728244966
Rh002_012_007+    hidden_activ_out_h001_012    tia_h_in_002_007+    14891.053514611822
Rh002_012_007-    hidden_activ_out_h001_012    tia_h_in_002_007-    11803.540284178429
Rh002_013_007+    hidden_activ_out_h001_013    tia_h_in_002_007+    15125.370970914835
Rh002_013_007-    hidden_activ_out_h001_013    tia_h_in_002_007-    8068.622722995875
Rh002_014_007+    hidden_activ_out_h001_014    tia_h_in_002_007+    13402.653045394502
Rh002_014_007-    hidden_activ_out_h001_014    tia_h_in_002_007-    15096.876203976928
Rh002_015_007+    hidden_activ_out_h001_015    tia_h_in_002_007+    14939.013712170765
Rh002_015_007-    hidden_activ_out_h001_015    tia_h_in_002_007-    13034.228679242671
Rh002_016_007+    hidden_activ_out_h001_016    tia_h_in_002_007+    11020.538793623165
Rh002_016_007-    hidden_activ_out_h001_016    tia_h_in_002_007-    15000
Rh002_017_007+    hidden_activ_out_h001_017    tia_h_in_002_007+    14591.218169553977
Rh002_017_007-    hidden_activ_out_h001_017    tia_h_in_002_007-    15012.541905823684
Rh002_018_007+    hidden_activ_out_h001_018    tia_h_in_002_007+    15192.060304432298
Rh002_018_007-    hidden_activ_out_h001_018    tia_h_in_002_007-    11349.575138274231
Rh002_019_007+    hidden_activ_out_h001_019    tia_h_in_002_007+    10497.37046011438
Rh002_019_007-    hidden_activ_out_h001_019    tia_h_in_002_007-    15129.47460793589
Rh002_020_007+    hidden_activ_out_h001_020    tia_h_in_002_007+    15000
Rh002_020_007-    hidden_activ_out_h001_020    tia_h_in_002_007-    13467.43476967095

* Neuron 8
Rh002_001_008+    hidden_activ_out_h001_001    tia_h_in_002_008+    14488.322692703874
Rh002_001_008-    hidden_activ_out_h001_001    tia_h_in_002_008-    14935.170056093082
Rh002_002_008+    hidden_activ_out_h001_002    tia_h_in_002_008+    15071.065825206093
Rh002_002_008-    hidden_activ_out_h001_002    tia_h_in_002_008-    5435.983874341784
Rh002_003_008+    hidden_activ_out_h001_003    tia_h_in_002_008+    11142.866209793172
Rh002_003_008-    hidden_activ_out_h001_003    tia_h_in_002_008-    15018.95346269893
Rh002_004_008+    hidden_activ_out_h001_004    tia_h_in_002_008+    14102.100376665416
Rh002_004_008-    hidden_activ_out_h001_004    tia_h_in_002_008-    14865.411927602461
Rh002_005_008+    hidden_activ_out_h001_005    tia_h_in_002_008+    14927.371311304141
Rh002_005_008-    hidden_activ_out_h001_005    tia_h_in_002_008-    8354.539443515578
Rh002_006_008+    hidden_activ_out_h001_006    tia_h_in_002_008+    15045.165578073866
Rh002_006_008-    hidden_activ_out_h001_006    tia_h_in_002_008-    14115.564327018641
Rh002_007_008+    hidden_activ_out_h001_007    tia_h_in_002_008+    15152.967594935048
Rh002_007_008-    hidden_activ_out_h001_007    tia_h_in_002_008-    7355.315884754804
Rh002_008_008+    hidden_activ_out_h001_008    tia_h_in_002_008+    14810.201393031515
Rh002_008_008-    hidden_activ_out_h001_008    tia_h_in_002_008-    8320.149684905688
Rh002_009_008+    hidden_activ_out_h001_009    tia_h_in_002_008+    15305.610470704323
Rh002_009_008-    hidden_activ_out_h001_009    tia_h_in_002_008-    6295.052765603327
Rh002_010_008+    hidden_activ_out_h001_010    tia_h_in_002_008+    12790.063581958793
Rh002_010_008-    hidden_activ_out_h001_010    tia_h_in_002_008-    14980.334236388422
Rh002_011_008+    hidden_activ_out_h001_011    tia_h_in_002_008+    15070.892486562743
Rh002_011_008-    hidden_activ_out_h001_011    tia_h_in_002_008-    8262.163414024344
Rh002_012_008+    hidden_activ_out_h001_012    tia_h_in_002_008+    14992.345437880938
Rh002_012_008-    hidden_activ_out_h001_012    tia_h_in_002_008-    8216.070901333365
Rh002_013_008+    hidden_activ_out_h001_013    tia_h_in_002_008+    14942.10317757554
Rh002_013_008-    hidden_activ_out_h001_013    tia_h_in_002_008-    7082.180539944266
Rh002_014_008+    hidden_activ_out_h001_014    tia_h_in_002_008+    14001.61939586332
Rh002_014_008-    hidden_activ_out_h001_014    tia_h_in_002_008-    15083.945530556619
Rh002_015_008+    hidden_activ_out_h001_015    tia_h_in_002_008+    13098.01983617545
Rh002_015_008-    hidden_activ_out_h001_015    tia_h_in_002_008-    15149.279616243812
Rh002_016_008+    hidden_activ_out_h001_016    tia_h_in_002_008+    14996.744556448259
Rh002_016_008-    hidden_activ_out_h001_016    tia_h_in_002_008-    14697.23588782777
Rh002_017_008+    hidden_activ_out_h001_017    tia_h_in_002_008+    14981.539460242866
Rh002_017_008-    hidden_activ_out_h001_017    tia_h_in_002_008-    11949.558702392176
Rh002_018_008+    hidden_activ_out_h001_018    tia_h_in_002_008+    14853.196410289043
Rh002_018_008-    hidden_activ_out_h001_018    tia_h_in_002_008-    5914.832035321593
Rh002_019_008+    hidden_activ_out_h001_019    tia_h_in_002_008+    11388.227272750346
Rh002_019_008-    hidden_activ_out_h001_019    tia_h_in_002_008-    15000
Rh002_020_008+    hidden_activ_out_h001_020    tia_h_in_002_008+    15052.490390865107
Rh002_020_008-    hidden_activ_out_h001_020    tia_h_in_002_008-    6331.644532038367

* Neuron 9
Rh002_001_009+    hidden_activ_out_h001_001    tia_h_in_002_009+    14967.308085519697
Rh002_001_009-    hidden_activ_out_h001_001    tia_h_in_002_009-    14979.386495286619
Rh002_002_009+    hidden_activ_out_h001_002    tia_h_in_002_009+    15025.909559851365
Rh002_002_009-    hidden_activ_out_h001_002    tia_h_in_002_009-    6934.129875476963
Rh002_003_009+    hidden_activ_out_h001_003    tia_h_in_002_009+    9795.901351869294
Rh002_003_009-    hidden_activ_out_h001_003    tia_h_in_002_009-    15190.940055179597
Rh002_004_009+    hidden_activ_out_h001_004    tia_h_in_002_009+    15050.855758376905
Rh002_004_009-    hidden_activ_out_h001_004    tia_h_in_002_009-    14406.29738907017
Rh002_005_009+    hidden_activ_out_h001_005    tia_h_in_002_009+    14990.828744489056
Rh002_005_009-    hidden_activ_out_h001_005    tia_h_in_002_009-    7602.349930282262
Rh002_006_009+    hidden_activ_out_h001_006    tia_h_in_002_009+    12991.266263165742
Rh002_006_009-    hidden_activ_out_h001_006    tia_h_in_002_009-    14992.666670771487
Rh002_007_009+    hidden_activ_out_h001_007    tia_h_in_002_009+    14955.004319514008
Rh002_007_009-    hidden_activ_out_h001_007    tia_h_in_002_009-    8502.26547460122
Rh002_008_009+    hidden_activ_out_h001_008    tia_h_in_002_009+    5000
Rh002_008_009-    hidden_activ_out_h001_008    tia_h_in_002_009-    8618.608273907525
Rh002_009_009+    hidden_activ_out_h001_009    tia_h_in_002_009+    15054.72974661448
Rh002_009_009-    hidden_activ_out_h001_009    tia_h_in_002_009-    7219.335949814323
Rh002_010_009+    hidden_activ_out_h001_010    tia_h_in_002_009+    13352.918701430366
Rh002_010_009-    hidden_activ_out_h001_010    tia_h_in_002_009-    15051.008170626383
Rh002_011_009+    hidden_activ_out_h001_011    tia_h_in_002_009+    15000
Rh002_011_009-    hidden_activ_out_h001_011    tia_h_in_002_009-    8001.133140847763
Rh002_012_009+    hidden_activ_out_h001_012    tia_h_in_002_009+    5000
Rh002_012_009-    hidden_activ_out_h001_012    tia_h_in_002_009-    5000
Rh002_013_009+    hidden_activ_out_h001_013    tia_h_in_002_009+    15087.750695512445
Rh002_013_009-    hidden_activ_out_h001_013    tia_h_in_002_009-    6733.421768182898
Rh002_014_009+    hidden_activ_out_h001_014    tia_h_in_002_009+    13749.692142024966
Rh002_014_009-    hidden_activ_out_h001_014    tia_h_in_002_009-    15055.215685897121
Rh002_015_009+    hidden_activ_out_h001_015    tia_h_in_002_009+    15081.841048562479
Rh002_015_009-    hidden_activ_out_h001_015    tia_h_in_002_009-    14867.137293847107
Rh002_016_009+    hidden_activ_out_h001_016    tia_h_in_002_009+    15178.111930303286
Rh002_016_009-    hidden_activ_out_h001_016    tia_h_in_002_009-    15000
Rh002_017_009+    hidden_activ_out_h001_017    tia_h_in_002_009+    15081.548022136585
Rh002_017_009-    hidden_activ_out_h001_017    tia_h_in_002_009-    14848.550278419463
Rh002_018_009+    hidden_activ_out_h001_018    tia_h_in_002_009+    14811.822029612229
Rh002_018_009-    hidden_activ_out_h001_018    tia_h_in_002_009-    8907.886533822983
Rh002_019_009+    hidden_activ_out_h001_019    tia_h_in_002_009+    11277.805867632931
Rh002_019_009-    hidden_activ_out_h001_019    tia_h_in_002_009-    15014.449186606582
Rh002_020_009+    hidden_activ_out_h001_020    tia_h_in_002_009+    14928.383269039134
Rh002_020_009-    hidden_activ_out_h001_020    tia_h_in_002_009-    11910.655816822573

* Neuron 10
Rh002_001_010+    hidden_activ_out_h001_001    tia_h_in_002_010+    9039.658974211798
Rh002_001_010-    hidden_activ_out_h001_001    tia_h_in_002_010-    14885.758042319567
Rh002_002_010+    hidden_activ_out_h001_002    tia_h_in_002_010+    14921.340263540613
Rh002_002_010-    hidden_activ_out_h001_002    tia_h_in_002_010-    5000
Rh002_003_010+    hidden_activ_out_h001_003    tia_h_in_002_010+    10373.781090957527
Rh002_003_010-    hidden_activ_out_h001_003    tia_h_in_002_010-    15065.782239219821
Rh002_004_010+    hidden_activ_out_h001_004    tia_h_in_002_010+    13345.075413146753
Rh002_004_010-    hidden_activ_out_h001_004    tia_h_in_002_010-    5000
Rh002_005_010+    hidden_activ_out_h001_005    tia_h_in_002_010+    14945.476296284924
Rh002_005_010-    hidden_activ_out_h001_005    tia_h_in_002_010-    9178.782968237714
Rh002_006_010+    hidden_activ_out_h001_006    tia_h_in_002_010+    12872.08694170224
Rh002_006_010-    hidden_activ_out_h001_006    tia_h_in_002_010-    15126.176826050001
Rh002_007_010+    hidden_activ_out_h001_007    tia_h_in_002_010+    14995.235375270931
Rh002_007_010-    hidden_activ_out_h001_007    tia_h_in_002_010-    11147.713890046722
Rh002_008_010+    hidden_activ_out_h001_008    tia_h_in_002_010+    14925.172569154282
Rh002_008_010-    hidden_activ_out_h001_008    tia_h_in_002_010-    9995.406817529014
Rh002_009_010+    hidden_activ_out_h001_009    tia_h_in_002_010+    15120.489927134735
Rh002_009_010-    hidden_activ_out_h001_009    tia_h_in_002_010-    12715.209651513025
Rh002_010_010+    hidden_activ_out_h001_010    tia_h_in_002_010+    15021.571539873994
Rh002_010_010-    hidden_activ_out_h001_010    tia_h_in_002_010-    13346.089310383913
Rh002_011_010+    hidden_activ_out_h001_011    tia_h_in_002_010+    15066.40611674338
Rh002_011_010-    hidden_activ_out_h001_011    tia_h_in_002_010-    11339.778206807729
Rh002_012_010+    hidden_activ_out_h001_012    tia_h_in_002_010+    14959.763852930355
Rh002_012_010-    hidden_activ_out_h001_012    tia_h_in_002_010-    14186.396769014202
Rh002_013_010+    hidden_activ_out_h001_013    tia_h_in_002_010+    14915.93267529797
Rh002_013_010-    hidden_activ_out_h001_013    tia_h_in_002_010-    11909.105138495075
Rh002_014_010+    hidden_activ_out_h001_014    tia_h_in_002_010+    14554.530014882825
Rh002_014_010-    hidden_activ_out_h001_014    tia_h_in_002_010-    5000
Rh002_015_010+    hidden_activ_out_h001_015    tia_h_in_002_010+    13388.37568627647
Rh002_015_010-    hidden_activ_out_h001_015    tia_h_in_002_010-    14926.669832163008
Rh002_016_010+    hidden_activ_out_h001_016    tia_h_in_002_010+    9012.29610021588
Rh002_016_010-    hidden_activ_out_h001_016    tia_h_in_002_010-    15314.769151592689
Rh002_017_010+    hidden_activ_out_h001_017    tia_h_in_002_010+    10753.910950276997
Rh002_017_010-    hidden_activ_out_h001_017    tia_h_in_002_010-    14776.360995751353
Rh002_018_010+    hidden_activ_out_h001_018    tia_h_in_002_010+    15003.655781910058
Rh002_018_010-    hidden_activ_out_h001_018    tia_h_in_002_010-    14099.21288766676
Rh002_019_010+    hidden_activ_out_h001_019    tia_h_in_002_010+    5000
Rh002_019_010-    hidden_activ_out_h001_019    tia_h_in_002_010-    5000
Rh002_020_010+    hidden_activ_out_h001_020    tia_h_in_002_010+    14913.249049831178
Rh002_020_010-    hidden_activ_out_h001_020    tia_h_in_002_010-    5000

* ----- Bias
    
        
Rb_h002_001+    b_002    tia_h_in_002_001+    12907.992158871493
Rb_h002_001-    b_002    tia_h_in_002_001-    15049.026920717279
Rb_h002_002+    b_002    tia_h_in_002_002+    12276.76559975711
Rb_h002_002-    b_002    tia_h_in_002_002-    15091.634744561383
Rb_h002_003+    b_002    tia_h_in_002_003+    12277.58140996887
Rb_h002_003-    b_002    tia_h_in_002_003-    15022.29035466802
Rb_h002_004+    b_002    tia_h_in_002_004+    13960.006055339856
Rb_h002_004-    b_002    tia_h_in_002_004-    14877.370133635255
Rb_h002_005+    b_002    tia_h_in_002_005+    13960.566771213287
Rb_h002_005-    b_002    tia_h_in_002_005-    15024.270351927595
Rb_h002_006+    b_002    tia_h_in_002_006+    13200.904218689844
Rb_h002_006-    b_002    tia_h_in_002_006-    15033.441590185848
Rb_h002_007+    b_002    tia_h_in_002_007+    12012.84927883461
Rb_h002_007-    b_002    tia_h_in_002_007-    14965.755893392816
Rb_h002_008+    b_002    tia_h_in_002_008+    11426.441680037584
Rb_h002_008-    b_002    tia_h_in_002_008-    15147.322502808078
Rb_h002_009+    b_002    tia_h_in_002_009+    11718.48707508234
Rb_h002_009-    b_002    tia_h_in_002_009-    14913.463109421427
Rb_h002_010+    b_002    tia_h_in_002_010+    13739.98098555697
Rb_h002_010-    b_002    tia_h_in_002_010-    15091.183320951488

* ----- Weights
* Layer 003

* Neuron 1
Rh003_001_001+    hidden_activ_out_h002_001    tia_h_in_003_001+    5000
Rh003_001_001-    hidden_activ_out_h002_001    tia_h_in_003_001-    5605.142949373137
Rh003_002_001+    hidden_activ_out_h002_002    tia_h_in_003_001+    4983.723487476977
Rh003_002_001-    hidden_activ_out_h002_002    tia_h_in_003_001-    15031.527355344855
Rh003_003_001+    hidden_activ_out_h002_003    tia_h_in_003_001+    15000
Rh003_003_001-    hidden_activ_out_h002_003    tia_h_in_003_001-    14800.491125088198
Rh003_004_001+    hidden_activ_out_h002_004    tia_h_in_003_001+    9118.899900040566
Rh003_004_001-    hidden_activ_out_h002_004    tia_h_in_003_001-    15000
Rh003_005_001+    hidden_activ_out_h002_005    tia_h_in_003_001+    8142.2079768851
Rh003_005_001-    hidden_activ_out_h002_005    tia_h_in_003_001-    15155.759009078862
Rh003_006_001+    hidden_activ_out_h002_006    tia_h_in_003_001+    14945.461104777813
Rh003_006_001-    hidden_activ_out_h002_006    tia_h_in_003_001-    5519.747174229925
Rh003_007_001+    hidden_activ_out_h002_007    tia_h_in_003_001+    7383.82099211443
Rh003_007_001-    hidden_activ_out_h002_007    tia_h_in_003_001-    14778.899477932344
Rh003_008_001+    hidden_activ_out_h002_008    tia_h_in_003_001+    5711.286898724222
Rh003_008_001-    hidden_activ_out_h002_008    tia_h_in_003_001-    15003.641295169644
Rh003_009_001+    hidden_activ_out_h002_009    tia_h_in_003_001+    6341.114397133808
Rh003_009_001-    hidden_activ_out_h002_009    tia_h_in_003_001-    15034.545134387865
Rh003_010_001+    hidden_activ_out_h002_010    tia_h_in_003_001+    8571.465492159547
Rh003_010_001-    hidden_activ_out_h002_010    tia_h_in_003_001-    15011.637082896574

* ----- Bias
    
        
Rb_h003_001+    b_003    tia_h_in_003_001+    14814.04023569448
Rb_h003_001-    b_003    tia_h_in_003_001-    6586.099692657345


* ----- Difference (V(R+) - V(R-))

* Layer 000
* Neuron 1
Rh001_fb_001+     tia_h_in_001_001+ tia_h_out_001_001+ 6000
Rh001_fb_001-     tia_h_in_001_001- tia_h_out_001_001- 6000
XUh001_001+       0 tia_h_in_001_001+ Vcc+ Vcc- tia_h_out_001_001+ Ve OPA684_0
XUh001_001-       0 tia_h_in_001_001- Vcc+ Vcc- tia_h_out_001_001- Ve OPA684_0
Rh001_sum_001+    tia_h_out_001_001+ sum_h_in_001_001- 260
Rh001_sum_001-    tia_h_out_001_001- sum_h_in_001_001+ 260
Rh001_sum_l_001   sum_h_in_001_001+ 0 745.2156186103822
Rh001_sum_fb_001  sum_h_in_001_001- sum_h_out_001_001 745.2156186103822
XUh001_sum_001    sum_h_in_001_001+ sum_h_in_001_001- Vcc+ Vcc- sum_h_out_001_001 MAX4223
* Neuron 2
Rh001_fb_002+     tia_h_in_001_002+ tia_h_out_001_002+ 6000
Rh001_fb_002-     tia_h_in_001_002- tia_h_out_001_002- 6000
XUh001_002+       0 tia_h_in_001_002+ Vcc+ Vcc- tia_h_out_001_002+ Ve OPA684_0
XUh001_002-       0 tia_h_in_001_002- Vcc+ Vcc- tia_h_out_001_002- Ve OPA684_0
Rh001_sum_002+    tia_h_out_001_002+ sum_h_in_001_002- 260
Rh001_sum_002-    tia_h_out_001_002- sum_h_in_001_002+ 260
Rh001_sum_l_002   sum_h_in_001_002+ 0 745.2156186103822
Rh001_sum_fb_002  sum_h_in_001_002- sum_h_out_001_002 745.2156186103822
XUh001_sum_002    sum_h_in_001_002+ sum_h_in_001_002- Vcc+ Vcc- sum_h_out_001_002 MAX4223
* Neuron 3
Rh001_fb_003+     tia_h_in_001_003+ tia_h_out_001_003+ 6000
Rh001_fb_003-     tia_h_in_001_003- tia_h_out_001_003- 6000
XUh001_003+       0 tia_h_in_001_003+ Vcc+ Vcc- tia_h_out_001_003+ Ve OPA684_0
XUh001_003-       0 tia_h_in_001_003- Vcc+ Vcc- tia_h_out_001_003- Ve OPA684_0
Rh001_sum_003+    tia_h_out_001_003+ sum_h_in_001_003- 260
Rh001_sum_003-    tia_h_out_001_003- sum_h_in_001_003+ 260
Rh001_sum_l_003   sum_h_in_001_003+ 0 745.2156186103822
Rh001_sum_fb_003  sum_h_in_001_003- sum_h_out_001_003 745.2156186103822
XUh001_sum_003    sum_h_in_001_003+ sum_h_in_001_003- Vcc+ Vcc- sum_h_out_001_003 MAX4223
* Neuron 4
Rh001_fb_004+     tia_h_in_001_004+ tia_h_out_001_004+ 6000
Rh001_fb_004-     tia_h_in_001_004- tia_h_out_001_004- 6000
XUh001_004+       0 tia_h_in_001_004+ Vcc+ Vcc- tia_h_out_001_004+ Ve OPA684_0
XUh001_004-       0 tia_h_in_001_004- Vcc+ Vcc- tia_h_out_001_004- Ve OPA684_0
Rh001_sum_004+    tia_h_out_001_004+ sum_h_in_001_004- 260
Rh001_sum_004-    tia_h_out_001_004- sum_h_in_001_004+ 260
Rh001_sum_l_004   sum_h_in_001_004+ 0 745.2156186103822
Rh001_sum_fb_004  sum_h_in_001_004- sum_h_out_001_004 745.2156186103822
XUh001_sum_004    sum_h_in_001_004+ sum_h_in_001_004- Vcc+ Vcc- sum_h_out_001_004 MAX4223
* Neuron 5
Rh001_fb_005+     tia_h_in_001_005+ tia_h_out_001_005+ 6000
Rh001_fb_005-     tia_h_in_001_005- tia_h_out_001_005- 6000
XUh001_005+       0 tia_h_in_001_005+ Vcc+ Vcc- tia_h_out_001_005+ Ve OPA684_0
XUh001_005-       0 tia_h_in_001_005- Vcc+ Vcc- tia_h_out_001_005- Ve OPA684_0
Rh001_sum_005+    tia_h_out_001_005+ sum_h_in_001_005- 260
Rh001_sum_005-    tia_h_out_001_005- sum_h_in_001_005+ 260
Rh001_sum_l_005   sum_h_in_001_005+ 0 745.2156186103822
Rh001_sum_fb_005  sum_h_in_001_005- sum_h_out_001_005 745.2156186103822
XUh001_sum_005    sum_h_in_001_005+ sum_h_in_001_005- Vcc+ Vcc- sum_h_out_001_005 MAX4223
* Neuron 6
Rh001_fb_006+     tia_h_in_001_006+ tia_h_out_001_006+ 6000
Rh001_fb_006-     tia_h_in_001_006- tia_h_out_001_006- 6000
XUh001_006+       0 tia_h_in_001_006+ Vcc+ Vcc- tia_h_out_001_006+ Ve OPA684_0
XUh001_006-       0 tia_h_in_001_006- Vcc+ Vcc- tia_h_out_001_006- Ve OPA684_0
Rh001_sum_006+    tia_h_out_001_006+ sum_h_in_001_006- 260
Rh001_sum_006-    tia_h_out_001_006- sum_h_in_001_006+ 260
Rh001_sum_l_006   sum_h_in_001_006+ 0 745.2156186103822
Rh001_sum_fb_006  sum_h_in_001_006- sum_h_out_001_006 745.2156186103822
XUh001_sum_006    sum_h_in_001_006+ sum_h_in_001_006- Vcc+ Vcc- sum_h_out_001_006 MAX4223
* Neuron 7
Rh001_fb_007+     tia_h_in_001_007+ tia_h_out_001_007+ 6000
Rh001_fb_007-     tia_h_in_001_007- tia_h_out_001_007- 6000
XUh001_007+       0 tia_h_in_001_007+ Vcc+ Vcc- tia_h_out_001_007+ Ve OPA684_0
XUh001_007-       0 tia_h_in_001_007- Vcc+ Vcc- tia_h_out_001_007- Ve OPA684_0
Rh001_sum_007+    tia_h_out_001_007+ sum_h_in_001_007- 260
Rh001_sum_007-    tia_h_out_001_007- sum_h_in_001_007+ 260
Rh001_sum_l_007   sum_h_in_001_007+ 0 745.2156186103822
Rh001_sum_fb_007  sum_h_in_001_007- sum_h_out_001_007 745.2156186103822
XUh001_sum_007    sum_h_in_001_007+ sum_h_in_001_007- Vcc+ Vcc- sum_h_out_001_007 MAX4223
* Neuron 8
Rh001_fb_008+     tia_h_in_001_008+ tia_h_out_001_008+ 6000
Rh001_fb_008-     tia_h_in_001_008- tia_h_out_001_008- 6000
XUh001_008+       0 tia_h_in_001_008+ Vcc+ Vcc- tia_h_out_001_008+ Ve OPA684_0
XUh001_008-       0 tia_h_in_001_008- Vcc+ Vcc- tia_h_out_001_008- Ve OPA684_0
Rh001_sum_008+    tia_h_out_001_008+ sum_h_in_001_008- 260
Rh001_sum_008-    tia_h_out_001_008- sum_h_in_001_008+ 260
Rh001_sum_l_008   sum_h_in_001_008+ 0 745.2156186103822
Rh001_sum_fb_008  sum_h_in_001_008- sum_h_out_001_008 745.2156186103822
XUh001_sum_008    sum_h_in_001_008+ sum_h_in_001_008- Vcc+ Vcc- sum_h_out_001_008 MAX4223
* Neuron 9
Rh001_fb_009+     tia_h_in_001_009+ tia_h_out_001_009+ 6000
Rh001_fb_009-     tia_h_in_001_009- tia_h_out_001_009- 6000
XUh001_009+       0 tia_h_in_001_009+ Vcc+ Vcc- tia_h_out_001_009+ Ve OPA684_0
XUh001_009-       0 tia_h_in_001_009- Vcc+ Vcc- tia_h_out_001_009- Ve OPA684_0
Rh001_sum_009+    tia_h_out_001_009+ sum_h_in_001_009- 260
Rh001_sum_009-    tia_h_out_001_009- sum_h_in_001_009+ 260
Rh001_sum_l_009   sum_h_in_001_009+ 0 745.2156186103822
Rh001_sum_fb_009  sum_h_in_001_009- sum_h_out_001_009 745.2156186103822
XUh001_sum_009    sum_h_in_001_009+ sum_h_in_001_009- Vcc+ Vcc- sum_h_out_001_009 MAX4223
* Neuron 10
Rh001_fb_010+     tia_h_in_001_010+ tia_h_out_001_010+ 6000
Rh001_fb_010-     tia_h_in_001_010- tia_h_out_001_010- 6000
XUh001_010+       0 tia_h_in_001_010+ Vcc+ Vcc- tia_h_out_001_010+ Ve OPA684_0
XUh001_010-       0 tia_h_in_001_010- Vcc+ Vcc- tia_h_out_001_010- Ve OPA684_0
Rh001_sum_010+    tia_h_out_001_010+ sum_h_in_001_010- 260
Rh001_sum_010-    tia_h_out_001_010- sum_h_in_001_010+ 260
Rh001_sum_l_010   sum_h_in_001_010+ 0 745.2156186103822
Rh001_sum_fb_010  sum_h_in_001_010- sum_h_out_001_010 745.2156186103822
XUh001_sum_010    sum_h_in_001_010+ sum_h_in_001_010- Vcc+ Vcc- sum_h_out_001_010 MAX4223
* Neuron 11
Rh001_fb_011+     tia_h_in_001_011+ tia_h_out_001_011+ 6000
Rh001_fb_011-     tia_h_in_001_011- tia_h_out_001_011- 6000
XUh001_011+       0 tia_h_in_001_011+ Vcc+ Vcc- tia_h_out_001_011+ Ve OPA684_0
XUh001_011-       0 tia_h_in_001_011- Vcc+ Vcc- tia_h_out_001_011- Ve OPA684_0
Rh001_sum_011+    tia_h_out_001_011+ sum_h_in_001_011- 260
Rh001_sum_011-    tia_h_out_001_011- sum_h_in_001_011+ 260
Rh001_sum_l_011   sum_h_in_001_011+ 0 745.2156186103822
Rh001_sum_fb_011  sum_h_in_001_011- sum_h_out_001_011 745.2156186103822
XUh001_sum_011    sum_h_in_001_011+ sum_h_in_001_011- Vcc+ Vcc- sum_h_out_001_011 MAX4223
* Neuron 12
Rh001_fb_012+     tia_h_in_001_012+ tia_h_out_001_012+ 6000
Rh001_fb_012-     tia_h_in_001_012- tia_h_out_001_012- 6000
XUh001_012+       0 tia_h_in_001_012+ Vcc+ Vcc- tia_h_out_001_012+ Ve OPA684_0
XUh001_012-       0 tia_h_in_001_012- Vcc+ Vcc- tia_h_out_001_012- Ve OPA684_0
Rh001_sum_012+    tia_h_out_001_012+ sum_h_in_001_012- 260
Rh001_sum_012-    tia_h_out_001_012- sum_h_in_001_012+ 260
Rh001_sum_l_012   sum_h_in_001_012+ 0 745.2156186103822
Rh001_sum_fb_012  sum_h_in_001_012- sum_h_out_001_012 745.2156186103822
XUh001_sum_012    sum_h_in_001_012+ sum_h_in_001_012- Vcc+ Vcc- sum_h_out_001_012 MAX4223
* Neuron 13
Rh001_fb_013+     tia_h_in_001_013+ tia_h_out_001_013+ 6000
Rh001_fb_013-     tia_h_in_001_013- tia_h_out_001_013- 6000
XUh001_013+       0 tia_h_in_001_013+ Vcc+ Vcc- tia_h_out_001_013+ Ve OPA684_0
XUh001_013-       0 tia_h_in_001_013- Vcc+ Vcc- tia_h_out_001_013- Ve OPA684_0
Rh001_sum_013+    tia_h_out_001_013+ sum_h_in_001_013- 260
Rh001_sum_013-    tia_h_out_001_013- sum_h_in_001_013+ 260
Rh001_sum_l_013   sum_h_in_001_013+ 0 745.2156186103822
Rh001_sum_fb_013  sum_h_in_001_013- sum_h_out_001_013 745.2156186103822
XUh001_sum_013    sum_h_in_001_013+ sum_h_in_001_013- Vcc+ Vcc- sum_h_out_001_013 MAX4223
* Neuron 14
Rh001_fb_014+     tia_h_in_001_014+ tia_h_out_001_014+ 6000
Rh001_fb_014-     tia_h_in_001_014- tia_h_out_001_014- 6000
XUh001_014+       0 tia_h_in_001_014+ Vcc+ Vcc- tia_h_out_001_014+ Ve OPA684_0
XUh001_014-       0 tia_h_in_001_014- Vcc+ Vcc- tia_h_out_001_014- Ve OPA684_0
Rh001_sum_014+    tia_h_out_001_014+ sum_h_in_001_014- 260
Rh001_sum_014-    tia_h_out_001_014- sum_h_in_001_014+ 260
Rh001_sum_l_014   sum_h_in_001_014+ 0 745.2156186103822
Rh001_sum_fb_014  sum_h_in_001_014- sum_h_out_001_014 745.2156186103822
XUh001_sum_014    sum_h_in_001_014+ sum_h_in_001_014- Vcc+ Vcc- sum_h_out_001_014 MAX4223
* Neuron 15
Rh001_fb_015+     tia_h_in_001_015+ tia_h_out_001_015+ 6000
Rh001_fb_015-     tia_h_in_001_015- tia_h_out_001_015- 6000
XUh001_015+       0 tia_h_in_001_015+ Vcc+ Vcc- tia_h_out_001_015+ Ve OPA684_0
XUh001_015-       0 tia_h_in_001_015- Vcc+ Vcc- tia_h_out_001_015- Ve OPA684_0
Rh001_sum_015+    tia_h_out_001_015+ sum_h_in_001_015- 260
Rh001_sum_015-    tia_h_out_001_015- sum_h_in_001_015+ 260
Rh001_sum_l_015   sum_h_in_001_015+ 0 745.2156186103822
Rh001_sum_fb_015  sum_h_in_001_015- sum_h_out_001_015 745.2156186103822
XUh001_sum_015    sum_h_in_001_015+ sum_h_in_001_015- Vcc+ Vcc- sum_h_out_001_015 MAX4223
* Neuron 16
Rh001_fb_016+     tia_h_in_001_016+ tia_h_out_001_016+ 6000
Rh001_fb_016-     tia_h_in_001_016- tia_h_out_001_016- 6000
XUh001_016+       0 tia_h_in_001_016+ Vcc+ Vcc- tia_h_out_001_016+ Ve OPA684_0
XUh001_016-       0 tia_h_in_001_016- Vcc+ Vcc- tia_h_out_001_016- Ve OPA684_0
Rh001_sum_016+    tia_h_out_001_016+ sum_h_in_001_016- 260
Rh001_sum_016-    tia_h_out_001_016- sum_h_in_001_016+ 260
Rh001_sum_l_016   sum_h_in_001_016+ 0 745.2156186103822
Rh001_sum_fb_016  sum_h_in_001_016- sum_h_out_001_016 745.2156186103822
XUh001_sum_016    sum_h_in_001_016+ sum_h_in_001_016- Vcc+ Vcc- sum_h_out_001_016 MAX4223
* Neuron 17
Rh001_fb_017+     tia_h_in_001_017+ tia_h_out_001_017+ 6000
Rh001_fb_017-     tia_h_in_001_017- tia_h_out_001_017- 6000
XUh001_017+       0 tia_h_in_001_017+ Vcc+ Vcc- tia_h_out_001_017+ Ve OPA684_0
XUh001_017-       0 tia_h_in_001_017- Vcc+ Vcc- tia_h_out_001_017- Ve OPA684_0
Rh001_sum_017+    tia_h_out_001_017+ sum_h_in_001_017- 260
Rh001_sum_017-    tia_h_out_001_017- sum_h_in_001_017+ 260
Rh001_sum_l_017   sum_h_in_001_017+ 0 745.2156186103822
Rh001_sum_fb_017  sum_h_in_001_017- sum_h_out_001_017 745.2156186103822
XUh001_sum_017    sum_h_in_001_017+ sum_h_in_001_017- Vcc+ Vcc- sum_h_out_001_017 MAX4223
* Neuron 18
Rh001_fb_018+     tia_h_in_001_018+ tia_h_out_001_018+ 6000
Rh001_fb_018-     tia_h_in_001_018- tia_h_out_001_018- 6000
XUh001_018+       0 tia_h_in_001_018+ Vcc+ Vcc- tia_h_out_001_018+ Ve OPA684_0
XUh001_018-       0 tia_h_in_001_018- Vcc+ Vcc- tia_h_out_001_018- Ve OPA684_0
Rh001_sum_018+    tia_h_out_001_018+ sum_h_in_001_018- 260
Rh001_sum_018-    tia_h_out_001_018- sum_h_in_001_018+ 260
Rh001_sum_l_018   sum_h_in_001_018+ 0 745.2156186103822
Rh001_sum_fb_018  sum_h_in_001_018- sum_h_out_001_018 745.2156186103822
XUh001_sum_018    sum_h_in_001_018+ sum_h_in_001_018- Vcc+ Vcc- sum_h_out_001_018 MAX4223
* Neuron 19
Rh001_fb_019+     tia_h_in_001_019+ tia_h_out_001_019+ 6000
Rh001_fb_019-     tia_h_in_001_019- tia_h_out_001_019- 6000
XUh001_019+       0 tia_h_in_001_019+ Vcc+ Vcc- tia_h_out_001_019+ Ve OPA684_0
XUh001_019-       0 tia_h_in_001_019- Vcc+ Vcc- tia_h_out_001_019- Ve OPA684_0
Rh001_sum_019+    tia_h_out_001_019+ sum_h_in_001_019- 260
Rh001_sum_019-    tia_h_out_001_019- sum_h_in_001_019+ 260
Rh001_sum_l_019   sum_h_in_001_019+ 0 745.2156186103822
Rh001_sum_fb_019  sum_h_in_001_019- sum_h_out_001_019 745.2156186103822
XUh001_sum_019    sum_h_in_001_019+ sum_h_in_001_019- Vcc+ Vcc- sum_h_out_001_019 MAX4223
* Neuron 20
Rh001_fb_020+     tia_h_in_001_020+ tia_h_out_001_020+ 6000
Rh001_fb_020-     tia_h_in_001_020- tia_h_out_001_020- 6000
XUh001_020+       0 tia_h_in_001_020+ Vcc+ Vcc- tia_h_out_001_020+ Ve OPA684_0
XUh001_020-       0 tia_h_in_001_020- Vcc+ Vcc- tia_h_out_001_020- Ve OPA684_0
Rh001_sum_020+    tia_h_out_001_020+ sum_h_in_001_020- 260
Rh001_sum_020-    tia_h_out_001_020- sum_h_in_001_020+ 260
Rh001_sum_l_020   sum_h_in_001_020+ 0 745.2156186103822
Rh001_sum_fb_020  sum_h_in_001_020- sum_h_out_001_020 745.2156186103822
XUh001_sum_020    sum_h_in_001_020+ sum_h_in_001_020- Vcc+ Vcc- sum_h_out_001_020 MAX4223

* Layer 001
* Neuron 1
Rh002_fb_001+     tia_h_in_002_001+ tia_h_out_002_001+ 6000
Rh002_fb_001-     tia_h_in_002_001- tia_h_out_002_001- 6000
XUh002_001+       0 tia_h_in_002_001+ Vcc+ Vcc- tia_h_out_002_001+ Ve OPA684_0
XUh002_001-       0 tia_h_in_002_001- Vcc+ Vcc- tia_h_out_002_001- Ve OPA684_0
Rh002_sum_001+    tia_h_out_002_001+ sum_h_in_002_001- 260
Rh002_sum_001-    tia_h_out_002_001- sum_h_in_002_001+ 260
Rh002_sum_l_001   sum_h_in_002_001+ 0 745.2156186103822
Rh002_sum_fb_001  sum_h_in_002_001- sum_h_out_002_001 745.2156186103822
XUh002_sum_001    sum_h_in_002_001+ sum_h_in_002_001- Vcc+ Vcc- sum_h_out_002_001 MAX4223
* Neuron 2
Rh002_fb_002+     tia_h_in_002_002+ tia_h_out_002_002+ 6000
Rh002_fb_002-     tia_h_in_002_002- tia_h_out_002_002- 6000
XUh002_002+       0 tia_h_in_002_002+ Vcc+ Vcc- tia_h_out_002_002+ Ve OPA684_0
XUh002_002-       0 tia_h_in_002_002- Vcc+ Vcc- tia_h_out_002_002- Ve OPA684_0
Rh002_sum_002+    tia_h_out_002_002+ sum_h_in_002_002- 260
Rh002_sum_002-    tia_h_out_002_002- sum_h_in_002_002+ 260
Rh002_sum_l_002   sum_h_in_002_002+ 0 745.2156186103822
Rh002_sum_fb_002  sum_h_in_002_002- sum_h_out_002_002 745.2156186103822
XUh002_sum_002    sum_h_in_002_002+ sum_h_in_002_002- Vcc+ Vcc- sum_h_out_002_002 MAX4223
* Neuron 3
Rh002_fb_003+     tia_h_in_002_003+ tia_h_out_002_003+ 6000
Rh002_fb_003-     tia_h_in_002_003- tia_h_out_002_003- 6000
XUh002_003+       0 tia_h_in_002_003+ Vcc+ Vcc- tia_h_out_002_003+ Ve OPA684_0
XUh002_003-       0 tia_h_in_002_003- Vcc+ Vcc- tia_h_out_002_003- Ve OPA684_0
Rh002_sum_003+    tia_h_out_002_003+ sum_h_in_002_003- 260
Rh002_sum_003-    tia_h_out_002_003- sum_h_in_002_003+ 260
Rh002_sum_l_003   sum_h_in_002_003+ 0 745.2156186103822
Rh002_sum_fb_003  sum_h_in_002_003- sum_h_out_002_003 745.2156186103822
XUh002_sum_003    sum_h_in_002_003+ sum_h_in_002_003- Vcc+ Vcc- sum_h_out_002_003 MAX4223
* Neuron 4
Rh002_fb_004+     tia_h_in_002_004+ tia_h_out_002_004+ 6000
Rh002_fb_004-     tia_h_in_002_004- tia_h_out_002_004- 6000
XUh002_004+       0 tia_h_in_002_004+ Vcc+ Vcc- tia_h_out_002_004+ Ve OPA684_0
XUh002_004-       0 tia_h_in_002_004- Vcc+ Vcc- tia_h_out_002_004- Ve OPA684_0
Rh002_sum_004+    tia_h_out_002_004+ sum_h_in_002_004- 260
Rh002_sum_004-    tia_h_out_002_004- sum_h_in_002_004+ 260
Rh002_sum_l_004   sum_h_in_002_004+ 0 745.2156186103822
Rh002_sum_fb_004  sum_h_in_002_004- sum_h_out_002_004 745.2156186103822
XUh002_sum_004    sum_h_in_002_004+ sum_h_in_002_004- Vcc+ Vcc- sum_h_out_002_004 MAX4223
* Neuron 5
Rh002_fb_005+     tia_h_in_002_005+ tia_h_out_002_005+ 6000
Rh002_fb_005-     tia_h_in_002_005- tia_h_out_002_005- 6000
XUh002_005+       0 tia_h_in_002_005+ Vcc+ Vcc- tia_h_out_002_005+ Ve OPA684_0
XUh002_005-       0 tia_h_in_002_005- Vcc+ Vcc- tia_h_out_002_005- Ve OPA684_0
Rh002_sum_005+    tia_h_out_002_005+ sum_h_in_002_005- 260
Rh002_sum_005-    tia_h_out_002_005- sum_h_in_002_005+ 260
Rh002_sum_l_005   sum_h_in_002_005+ 0 745.2156186103822
Rh002_sum_fb_005  sum_h_in_002_005- sum_h_out_002_005 745.2156186103822
XUh002_sum_005    sum_h_in_002_005+ sum_h_in_002_005- Vcc+ Vcc- sum_h_out_002_005 MAX4223
* Neuron 6
Rh002_fb_006+     tia_h_in_002_006+ tia_h_out_002_006+ 6000
Rh002_fb_006-     tia_h_in_002_006- tia_h_out_002_006- 6000
XUh002_006+       0 tia_h_in_002_006+ Vcc+ Vcc- tia_h_out_002_006+ Ve OPA684_0
XUh002_006-       0 tia_h_in_002_006- Vcc+ Vcc- tia_h_out_002_006- Ve OPA684_0
Rh002_sum_006+    tia_h_out_002_006+ sum_h_in_002_006- 260
Rh002_sum_006-    tia_h_out_002_006- sum_h_in_002_006+ 260
Rh002_sum_l_006   sum_h_in_002_006+ 0 745.2156186103822
Rh002_sum_fb_006  sum_h_in_002_006- sum_h_out_002_006 745.2156186103822
XUh002_sum_006    sum_h_in_002_006+ sum_h_in_002_006- Vcc+ Vcc- sum_h_out_002_006 MAX4223
* Neuron 7
Rh002_fb_007+     tia_h_in_002_007+ tia_h_out_002_007+ 6000
Rh002_fb_007-     tia_h_in_002_007- tia_h_out_002_007- 6000
XUh002_007+       0 tia_h_in_002_007+ Vcc+ Vcc- tia_h_out_002_007+ Ve OPA684_0
XUh002_007-       0 tia_h_in_002_007- Vcc+ Vcc- tia_h_out_002_007- Ve OPA684_0
Rh002_sum_007+    tia_h_out_002_007+ sum_h_in_002_007- 260
Rh002_sum_007-    tia_h_out_002_007- sum_h_in_002_007+ 260
Rh002_sum_l_007   sum_h_in_002_007+ 0 745.2156186103822
Rh002_sum_fb_007  sum_h_in_002_007- sum_h_out_002_007 745.2156186103822
XUh002_sum_007    sum_h_in_002_007+ sum_h_in_002_007- Vcc+ Vcc- sum_h_out_002_007 MAX4223
* Neuron 8
Rh002_fb_008+     tia_h_in_002_008+ tia_h_out_002_008+ 6000
Rh002_fb_008-     tia_h_in_002_008- tia_h_out_002_008- 6000
XUh002_008+       0 tia_h_in_002_008+ Vcc+ Vcc- tia_h_out_002_008+ Ve OPA684_0
XUh002_008-       0 tia_h_in_002_008- Vcc+ Vcc- tia_h_out_002_008- Ve OPA684_0
Rh002_sum_008+    tia_h_out_002_008+ sum_h_in_002_008- 260
Rh002_sum_008-    tia_h_out_002_008- sum_h_in_002_008+ 260
Rh002_sum_l_008   sum_h_in_002_008+ 0 745.2156186103822
Rh002_sum_fb_008  sum_h_in_002_008- sum_h_out_002_008 745.2156186103822
XUh002_sum_008    sum_h_in_002_008+ sum_h_in_002_008- Vcc+ Vcc- sum_h_out_002_008 MAX4223
* Neuron 9
Rh002_fb_009+     tia_h_in_002_009+ tia_h_out_002_009+ 6000
Rh002_fb_009-     tia_h_in_002_009- tia_h_out_002_009- 6000
XUh002_009+       0 tia_h_in_002_009+ Vcc+ Vcc- tia_h_out_002_009+ Ve OPA684_0
XUh002_009-       0 tia_h_in_002_009- Vcc+ Vcc- tia_h_out_002_009- Ve OPA684_0
Rh002_sum_009+    tia_h_out_002_009+ sum_h_in_002_009- 260
Rh002_sum_009-    tia_h_out_002_009- sum_h_in_002_009+ 260
Rh002_sum_l_009   sum_h_in_002_009+ 0 745.2156186103822
Rh002_sum_fb_009  sum_h_in_002_009- sum_h_out_002_009 745.2156186103822
XUh002_sum_009    sum_h_in_002_009+ sum_h_in_002_009- Vcc+ Vcc- sum_h_out_002_009 MAX4223
* Neuron 10
Rh002_fb_010+     tia_h_in_002_010+ tia_h_out_002_010+ 6000
Rh002_fb_010-     tia_h_in_002_010- tia_h_out_002_010- 6000
XUh002_010+       0 tia_h_in_002_010+ Vcc+ Vcc- tia_h_out_002_010+ Ve OPA684_0
XUh002_010-       0 tia_h_in_002_010- Vcc+ Vcc- tia_h_out_002_010- Ve OPA684_0
Rh002_sum_010+    tia_h_out_002_010+ sum_h_in_002_010- 260
Rh002_sum_010-    tia_h_out_002_010- sum_h_in_002_010+ 260
Rh002_sum_l_010   sum_h_in_002_010+ 0 745.2156186103822
Rh002_sum_fb_010  sum_h_in_002_010- sum_h_out_002_010 745.2156186103822
XUh002_sum_010    sum_h_in_002_010+ sum_h_in_002_010- Vcc+ Vcc- sum_h_out_002_010 MAX4223

* Layer 002
* Neuron 1
Rh003_fb_001+     tia_h_in_003_001+ tia_h_out_003_001+ 6000
Rh003_fb_001-     tia_h_in_003_001- tia_h_out_003_001- 6000
XUh003_001+       0 tia_h_in_003_001+ Vcc+ Vcc- tia_h_out_003_001+ Ve OPA684_0
XUh003_001-       0 tia_h_in_003_001- Vcc+ Vcc- tia_h_out_003_001- Ve OPA684_0
Rh003_sum_001+    tia_h_out_003_001+ sum_h_in_003_001- 260
Rh003_sum_001-    tia_h_out_003_001- sum_h_in_003_001+ 260
Rh003_sum_l_001   sum_h_in_003_001+ 0 745.2156186103822
Rh003_sum_fb_001  sum_h_in_003_001- sum_h_out_003_001 745.2156186103822
XUh003_sum_001    sum_h_in_003_001+ sum_h_in_003_001- Vcc+ Vcc- sum_h_out_003_001 MAX4223


* ----- Activation function Hard-Tanh)


* Layer 000
* Neuron 1
* XHardTanh_h001_001 sum_h_out_001_001 hidden_activ_out_h001_001 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_001 sum_h_out_001_001 hidden_activ_out_h001_001 ReLU
*XSigmoid_001_001 sum_h_out_001_001 hidden_activ_out_h001_001 RNN_Sigmoid3_HA
* Neuron 2
* XHardTanh_h001_002 sum_h_out_001_002 hidden_activ_out_h001_002 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_002 sum_h_out_001_002 hidden_activ_out_h001_002 ReLU
*XSigmoid_001_002 sum_h_out_001_002 hidden_activ_out_h001_002 RNN_Sigmoid3_HA
* Neuron 3
* XHardTanh_h001_003 sum_h_out_001_003 hidden_activ_out_h001_003 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_003 sum_h_out_001_003 hidden_activ_out_h001_003 ReLU
*XSigmoid_001_003 sum_h_out_001_003 hidden_activ_out_h001_003 RNN_Sigmoid3_HA
* Neuron 4
* XHardTanh_h001_004 sum_h_out_001_004 hidden_activ_out_h001_004 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_004 sum_h_out_001_004 hidden_activ_out_h001_004 ReLU
*XSigmoid_001_004 sum_h_out_001_004 hidden_activ_out_h001_004 RNN_Sigmoid3_HA
* Neuron 5
* XHardTanh_h001_005 sum_h_out_001_005 hidden_activ_out_h001_005 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_005 sum_h_out_001_005 hidden_activ_out_h001_005 ReLU
*XSigmoid_001_005 sum_h_out_001_005 hidden_activ_out_h001_005 RNN_Sigmoid3_HA
* Neuron 6
* XHardTanh_h001_006 sum_h_out_001_006 hidden_activ_out_h001_006 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_006 sum_h_out_001_006 hidden_activ_out_h001_006 ReLU
*XSigmoid_001_006 sum_h_out_001_006 hidden_activ_out_h001_006 RNN_Sigmoid3_HA
* Neuron 7
* XHardTanh_h001_007 sum_h_out_001_007 hidden_activ_out_h001_007 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_007 sum_h_out_001_007 hidden_activ_out_h001_007 ReLU
*XSigmoid_001_007 sum_h_out_001_007 hidden_activ_out_h001_007 RNN_Sigmoid3_HA
* Neuron 8
* XHardTanh_h001_008 sum_h_out_001_008 hidden_activ_out_h001_008 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_008 sum_h_out_001_008 hidden_activ_out_h001_008 ReLU
*XSigmoid_001_008 sum_h_out_001_008 hidden_activ_out_h001_008 RNN_Sigmoid3_HA
* Neuron 9
* XHardTanh_h001_009 sum_h_out_001_009 hidden_activ_out_h001_009 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_009 sum_h_out_001_009 hidden_activ_out_h001_009 ReLU
*XSigmoid_001_009 sum_h_out_001_009 hidden_activ_out_h001_009 RNN_Sigmoid3_HA
* Neuron 10
* XHardTanh_h001_010 sum_h_out_001_010 hidden_activ_out_h001_010 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_010 sum_h_out_001_010 hidden_activ_out_h001_010 ReLU
*XSigmoid_001_010 sum_h_out_001_010 hidden_activ_out_h001_010 RNN_Sigmoid3_HA
* Neuron 11
* XHardTanh_h001_011 sum_h_out_001_011 hidden_activ_out_h001_011 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_011 sum_h_out_001_011 hidden_activ_out_h001_011 ReLU
*XSigmoid_001_011 sum_h_out_001_011 hidden_activ_out_h001_011 RNN_Sigmoid3_HA
* Neuron 12
* XHardTanh_h001_012 sum_h_out_001_012 hidden_activ_out_h001_012 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_012 sum_h_out_001_012 hidden_activ_out_h001_012 ReLU
*XSigmoid_001_012 sum_h_out_001_012 hidden_activ_out_h001_012 RNN_Sigmoid3_HA
* Neuron 13
* XHardTanh_h001_013 sum_h_out_001_013 hidden_activ_out_h001_013 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_013 sum_h_out_001_013 hidden_activ_out_h001_013 ReLU
*XSigmoid_001_013 sum_h_out_001_013 hidden_activ_out_h001_013 RNN_Sigmoid3_HA
* Neuron 14
* XHardTanh_h001_014 sum_h_out_001_014 hidden_activ_out_h001_014 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_014 sum_h_out_001_014 hidden_activ_out_h001_014 ReLU
*XSigmoid_001_014 sum_h_out_001_014 hidden_activ_out_h001_014 RNN_Sigmoid3_HA
* Neuron 15
* XHardTanh_h001_015 sum_h_out_001_015 hidden_activ_out_h001_015 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_015 sum_h_out_001_015 hidden_activ_out_h001_015 ReLU
*XSigmoid_001_015 sum_h_out_001_015 hidden_activ_out_h001_015 RNN_Sigmoid3_HA
* Neuron 16
* XHardTanh_h001_016 sum_h_out_001_016 hidden_activ_out_h001_016 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_016 sum_h_out_001_016 hidden_activ_out_h001_016 ReLU
*XSigmoid_001_016 sum_h_out_001_016 hidden_activ_out_h001_016 RNN_Sigmoid3_HA
* Neuron 17
* XHardTanh_h001_017 sum_h_out_001_017 hidden_activ_out_h001_017 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_017 sum_h_out_001_017 hidden_activ_out_h001_017 ReLU
*XSigmoid_001_017 sum_h_out_001_017 hidden_activ_out_h001_017 RNN_Sigmoid3_HA
* Neuron 18
* XHardTanh_h001_018 sum_h_out_001_018 hidden_activ_out_h001_018 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_018 sum_h_out_001_018 hidden_activ_out_h001_018 ReLU
*XSigmoid_001_018 sum_h_out_001_018 hidden_activ_out_h001_018 RNN_Sigmoid3_HA
* Neuron 19
* XHardTanh_h001_019 sum_h_out_001_019 hidden_activ_out_h001_019 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_019 sum_h_out_001_019 hidden_activ_out_h001_019 ReLU
*XSigmoid_001_019 sum_h_out_001_019 hidden_activ_out_h001_019 RNN_Sigmoid3_HA
* Neuron 20
* XHardTanh_h001_020 sum_h_out_001_020 hidden_activ_out_h001_020 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_020 sum_h_out_001_020 hidden_activ_out_h001_020 ReLU
*XSigmoid_001_020 sum_h_out_001_020 hidden_activ_out_h001_020 RNN_Sigmoid3_HA

* Layer 001
* Neuron 1
* XHardTanh_h002_001 sum_h_out_002_001 hidden_activ_out_h002_001 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_001 sum_h_out_002_001 hidden_activ_out_h002_001 ReLU
*XSigmoid_002_001 sum_h_out_002_001 hidden_activ_out_h002_001 RNN_Sigmoid3_HA
* Neuron 2
* XHardTanh_h002_002 sum_h_out_002_002 hidden_activ_out_h002_002 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_002 sum_h_out_002_002 hidden_activ_out_h002_002 ReLU
*XSigmoid_002_002 sum_h_out_002_002 hidden_activ_out_h002_002 RNN_Sigmoid3_HA
* Neuron 3
* XHardTanh_h002_003 sum_h_out_002_003 hidden_activ_out_h002_003 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_003 sum_h_out_002_003 hidden_activ_out_h002_003 ReLU
*XSigmoid_002_003 sum_h_out_002_003 hidden_activ_out_h002_003 RNN_Sigmoid3_HA
* Neuron 4
* XHardTanh_h002_004 sum_h_out_002_004 hidden_activ_out_h002_004 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_004 sum_h_out_002_004 hidden_activ_out_h002_004 ReLU
*XSigmoid_002_004 sum_h_out_002_004 hidden_activ_out_h002_004 RNN_Sigmoid3_HA
* Neuron 5
* XHardTanh_h002_005 sum_h_out_002_005 hidden_activ_out_h002_005 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_005 sum_h_out_002_005 hidden_activ_out_h002_005 ReLU
*XSigmoid_002_005 sum_h_out_002_005 hidden_activ_out_h002_005 RNN_Sigmoid3_HA
* Neuron 6
* XHardTanh_h002_006 sum_h_out_002_006 hidden_activ_out_h002_006 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_006 sum_h_out_002_006 hidden_activ_out_h002_006 ReLU
*XSigmoid_002_006 sum_h_out_002_006 hidden_activ_out_h002_006 RNN_Sigmoid3_HA
* Neuron 7
* XHardTanh_h002_007 sum_h_out_002_007 hidden_activ_out_h002_007 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_007 sum_h_out_002_007 hidden_activ_out_h002_007 ReLU
*XSigmoid_002_007 sum_h_out_002_007 hidden_activ_out_h002_007 RNN_Sigmoid3_HA
* Neuron 8
* XHardTanh_h002_008 sum_h_out_002_008 hidden_activ_out_h002_008 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_008 sum_h_out_002_008 hidden_activ_out_h002_008 ReLU
*XSigmoid_002_008 sum_h_out_002_008 hidden_activ_out_h002_008 RNN_Sigmoid3_HA
* Neuron 9
* XHardTanh_h002_009 sum_h_out_002_009 hidden_activ_out_h002_009 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_009 sum_h_out_002_009 hidden_activ_out_h002_009 ReLU
*XSigmoid_002_009 sum_h_out_002_009 hidden_activ_out_h002_009 RNN_Sigmoid3_HA
* Neuron 10
* XHardTanh_h002_010 sum_h_out_002_010 hidden_activ_out_h002_010 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_010 sum_h_out_002_010 hidden_activ_out_h002_010 ReLU
*XSigmoid_002_010 sum_h_out_002_010 hidden_activ_out_h002_010 RNN_Sigmoid3_HA

* Layer 002
* Neuron 1
* XHardTanh_h003_001 sum_h_out_003_001 hidden_activ_out_h003_001 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_003_001 sum_h_out_003_001 hidden_activ_out_h003_001 ReLU
*XSigmoid_003_001 sum_h_out_003_001 hidden_activ_out_h003_001 RNN_Sigmoid3_HA


.END