* Netlist that describe the physical circuit (components and connexions between them) to simulate, in Xyce formalism.
* To make the translation from any network size, the circuit is scaled up automatically using Jinja template engine.
*
* Xyce: https://xyce.sandia.gov
* Jinja: https://jinja.palletsprojects.com

* ======================== Simulation parameters ==========================

.TRAN 0.30ns 331.00ns

* OPTIONS TIMEINT change the time integration parameters
* ERROPTION (If 0 Local Truncation Error is used)
* METHOD: Time integration method
* NLMIN, NLMAX:  lower and upper bound for the desired number of nonlinear iterations
* DELMAX: The maximum time step-size used
* This additional line allows to fix convergence problem but increases the simulation time
* List variables to save in the result table
.PRINT TRAN V(sum_h_out_003_001) V(hidden_activ_out_h003_001)
+ V(i_001) V(i_002) V(i_003) V(i_004) V(i_005) V(i_006) V(i_007) V(i_008) V(i_009) V(i_010) V(i_011) V(i_012) V(i_013) V(i_014) V(i_015) V(i_016) V(i_017) V(i_018) V(i_019) V(i_020) V(i_021) V(i_022) V(i_023) V(i_024) V(i_025) V(i_026) V(i_027) V(i_028) V(i_029) V(i_030) V(i_031) V(i_032) V(i_033) V(i_034) V(i_035) V(i_036) V(i_037) V(i_038) V(i_039) V(i_040) V(i_041) V(i_042) V(i_043) V(i_044) V(i_045) V(i_046) V(i_047) V(i_048) V(i_049) V(i_050) V(i_051) V(i_052) V(i_053) V(i_054) V(i_055) V(i_056) V(i_057) V(i_058) V(i_059) V(i_060) V(i_061) V(i_062) V(i_063) V(i_064)
+ V(sum_h_out_001_001) V(hidden_activ_out_h001_001) V(sum_h_out_001_002) V(hidden_activ_out_h001_002) V(sum_h_out_001_003) V(hidden_activ_out_h001_003) V(sum_h_out_001_004) V(hidden_activ_out_h001_004) V(sum_h_out_001_005) V(hidden_activ_out_h001_005) V(sum_h_out_001_006) V(hidden_activ_out_h001_006) V(sum_h_out_001_007) V(hidden_activ_out_h001_007) V(sum_h_out_001_008) V(hidden_activ_out_h001_008) V(sum_h_out_001_009) V(hidden_activ_out_h001_009) V(sum_h_out_001_010) V(hidden_activ_out_h001_010) V(sum_h_out_001_011) V(hidden_activ_out_h001_011) V(sum_h_out_001_012) V(hidden_activ_out_h001_012) V(sum_h_out_001_013) V(hidden_activ_out_h001_013) V(sum_h_out_001_014) V(hidden_activ_out_h001_014) V(sum_h_out_001_015) V(hidden_activ_out_h001_015) V(sum_h_out_001_016) V(hidden_activ_out_h001_016) V(sum_h_out_001_017) V(hidden_activ_out_h001_017) V(sum_h_out_001_018) V(hidden_activ_out_h001_018) V(sum_h_out_001_019) V(hidden_activ_out_h001_019) V(sum_h_out_001_020) V(hidden_activ_out_h001_020)
+ V(tia_h_out_001_001+) V(tia_h_out_001_001-) V(tia_h_out_001_002+) V(tia_h_out_001_002-) V(tia_h_out_001_003+) V(tia_h_out_001_003-) V(tia_h_out_001_004+) V(tia_h_out_001_004-) V(tia_h_out_001_005+) V(tia_h_out_001_005-) V(tia_h_out_001_006+) V(tia_h_out_001_006-) V(tia_h_out_001_007+) V(tia_h_out_001_007-) V(tia_h_out_001_008+) V(tia_h_out_001_008-) V(tia_h_out_001_009+) V(tia_h_out_001_009-) V(tia_h_out_001_010+) V(tia_h_out_001_010-) V(tia_h_out_001_011+) V(tia_h_out_001_011-) V(tia_h_out_001_012+) V(tia_h_out_001_012-) V(tia_h_out_001_013+) V(tia_h_out_001_013-) V(tia_h_out_001_014+) V(tia_h_out_001_014-) V(tia_h_out_001_015+) V(tia_h_out_001_015-) V(tia_h_out_001_016+) V(tia_h_out_001_016-) V(tia_h_out_001_017+) V(tia_h_out_001_017-) V(tia_h_out_001_018+) V(tia_h_out_001_018-) V(tia_h_out_001_019+) V(tia_h_out_001_019-) V(tia_h_out_001_020+) V(tia_h_out_001_020-)
+ V(b_001)
+ V(sum_h_out_002_001) V(hidden_activ_out_h002_001) V(sum_h_out_002_002) V(hidden_activ_out_h002_002) V(sum_h_out_002_003) V(hidden_activ_out_h002_003) V(sum_h_out_002_004) V(hidden_activ_out_h002_004) V(sum_h_out_002_005) V(hidden_activ_out_h002_005) V(sum_h_out_002_006) V(hidden_activ_out_h002_006) V(sum_h_out_002_007) V(hidden_activ_out_h002_007) V(sum_h_out_002_008) V(hidden_activ_out_h002_008) V(sum_h_out_002_009) V(hidden_activ_out_h002_009) V(sum_h_out_002_010) V(hidden_activ_out_h002_010)
+ V(tia_h_out_002_001+) V(tia_h_out_002_001-) V(tia_h_out_002_002+) V(tia_h_out_002_002-) V(tia_h_out_002_003+) V(tia_h_out_002_003-) V(tia_h_out_002_004+) V(tia_h_out_002_004-) V(tia_h_out_002_005+) V(tia_h_out_002_005-) V(tia_h_out_002_006+) V(tia_h_out_002_006-) V(tia_h_out_002_007+) V(tia_h_out_002_007-) V(tia_h_out_002_008+) V(tia_h_out_002_008-) V(tia_h_out_002_009+) V(tia_h_out_002_009-) V(tia_h_out_002_010+) V(tia_h_out_002_010-)
+ V(b_002)
+ V(sum_h_out_003_001) V(hidden_activ_out_h003_001)
+ V(tia_h_out_003_001+) V(tia_h_out_003_001-)
+ V(b_003)

* =============================== Models ==================================

* Call the defined components model from the specified path
*.INCLUDE "./components/MAX4223.sub"
.INCLUDE "./components/TLV3501.sub"
*.INCLUDE "./components/OPA684.sub"

* Import custom sub-circuits
.INCLUDE "./components/activations.sub"
.INCLUDE "./components/lumped_line.sub"
.INCLUDE "./components/Sigmoid3_HA.spice"

* Define diode model
.MODEL D_BAV74_1 D( IS=2.073F N=1 BV=50 IBV=100N RS=1.336 
+      CJO=2P VJ=750M M=330M FC=500M TT=5.771N 
+      EG=1.11 XTI=3 KF=0 AF=1 )

* ============================== Voltages =================================

* ----- Input pulses
* Vi_num: The input voltage as pulse sequences
Vi_001    i_001    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.067V 281.00ns 1.067V 301.00ns 1.050V 381.00ns 1.050V
Vi_002    i_002    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.062V 281.00ns 1.062V 301.00ns 1.050V 381.00ns 1.050V
Vi_003    i_003    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.134V 281.00ns 1.134V 301.00ns 1.050V 381.00ns 1.050V
Vi_004    i_004    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.119V 281.00ns 1.119V 301.00ns 1.050V 381.00ns 1.050V
Vi_005    i_005    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.205V 281.00ns 1.205V 301.00ns 1.050V 381.00ns 1.050V
Vi_006    i_006    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.181V 281.00ns 1.181V 301.00ns 1.050V 381.00ns 1.050V
Vi_007    i_007    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.177V 281.00ns 1.177V 301.00ns 1.050V 381.00ns 1.050V
Vi_008    i_008    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.225V 281.00ns 1.225V 301.00ns 1.050V 381.00ns 1.050V
Vi_009    i_009    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.058V 281.00ns 1.058V 301.00ns 1.050V 381.00ns 1.050V
Vi_010    i_010    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.062V 281.00ns 1.062V 301.00ns 1.050V 381.00ns 1.050V
Vi_011    i_011    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.136V 281.00ns 1.136V 301.00ns 1.050V 381.00ns 1.050V
Vi_012    i_012    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.113V 281.00ns 1.113V 301.00ns 1.050V 381.00ns 1.050V
Vi_013    i_013    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.211V 281.00ns 1.211V 301.00ns 1.050V 381.00ns 1.050V
Vi_014    i_014    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.175V 281.00ns 1.175V 301.00ns 1.050V 381.00ns 1.050V
Vi_015    i_015    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.157V 281.00ns 1.157V 301.00ns 1.050V 381.00ns 1.050V
Vi_016    i_016    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.238V 281.00ns 1.238V 301.00ns 1.050V 381.00ns 1.050V
Vi_017    i_017    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.064V 281.00ns 1.064V 301.00ns 1.050V 381.00ns 1.050V
Vi_018    i_018    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.126V 281.00ns 1.126V 301.00ns 1.050V 381.00ns 1.050V
Vi_019    i_019    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.092V 281.00ns 1.092V 301.00ns 1.050V 381.00ns 1.050V
Vi_020    i_020    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.119V 281.00ns 1.119V 301.00ns 1.050V 381.00ns 1.050V
Vi_021    i_021    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.201V 281.00ns 1.201V 301.00ns 1.050V 381.00ns 1.050V
Vi_022    i_022    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.139V 281.00ns 1.139V 301.00ns 1.050V 381.00ns 1.050V
Vi_023    i_023    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.113V 281.00ns 1.113V 301.00ns 1.050V 381.00ns 1.050V
Vi_024    i_024    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.278V 281.00ns 1.278V 301.00ns 1.050V 381.00ns 1.050V
Vi_025    i_025    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.050V 281.00ns 1.050V 301.00ns 1.050V 381.00ns 1.050V
Vi_026    i_026    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.146V 281.00ns 1.146V 301.00ns 1.050V 381.00ns 1.050V
Vi_027    i_027    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.135V 281.00ns 1.135V 301.00ns 1.050V 381.00ns 1.050V
Vi_028    i_028    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.162V 281.00ns 1.162V 301.00ns 1.050V 381.00ns 1.050V
Vi_029    i_029    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.212V 281.00ns 1.212V 301.00ns 1.050V 381.00ns 1.050V
Vi_030    i_030    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.178V 281.00ns 1.178V 301.00ns 1.050V 381.00ns 1.050V
Vi_031    i_031    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.149V 281.00ns 1.149V 301.00ns 1.050V 381.00ns 1.050V
Vi_032    i_032    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.296V 281.00ns 1.296V 301.00ns 1.050V 381.00ns 1.050V
Vi_033    i_033    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.063V 281.00ns 1.063V 301.00ns 1.050V 381.00ns 1.050V
Vi_034    i_034    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.135V 281.00ns 1.135V 301.00ns 1.050V 381.00ns 1.050V
Vi_035    i_035    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.129V 281.00ns 1.129V 301.00ns 1.050V 381.00ns 1.050V
Vi_036    i_036    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.202V 281.00ns 1.202V 301.00ns 1.050V 381.00ns 1.050V
Vi_037    i_037    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.252V 281.00ns 1.252V 301.00ns 1.050V 381.00ns 1.050V
Vi_038    i_038    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.208V 281.00ns 1.208V 301.00ns 1.050V 381.00ns 1.050V
Vi_039    i_039    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.138V 281.00ns 1.138V 301.00ns 1.050V 381.00ns 1.050V
Vi_040    i_040    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.295V 281.00ns 1.295V 301.00ns 1.050V 381.00ns 1.050V
Vi_041    i_041    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.108V 281.00ns 1.108V 301.00ns 1.050V 381.00ns 1.050V
Vi_042    i_042    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.128V 281.00ns 1.128V 301.00ns 1.050V 381.00ns 1.050V
Vi_043    i_043    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.144V 281.00ns 1.144V 301.00ns 1.050V 381.00ns 1.050V
Vi_044    i_044    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.200V 281.00ns 1.200V 301.00ns 1.050V 381.00ns 1.050V
Vi_045    i_045    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.257V 281.00ns 1.257V 301.00ns 1.050V 381.00ns 1.050V
Vi_046    i_046    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.199V 281.00ns 1.199V 301.00ns 1.050V 381.00ns 1.050V
Vi_047    i_047    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.220V 281.00ns 1.220V 301.00ns 1.050V 381.00ns 1.050V
Vi_048    i_048    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.298V 281.00ns 1.298V 301.00ns 1.050V 381.00ns 1.050V
Vi_049    i_049    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.102V 281.00ns 1.102V 301.00ns 1.050V 381.00ns 1.050V
Vi_050    i_050    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.115V 281.00ns 1.115V 301.00ns 1.050V 381.00ns 1.050V
Vi_051    i_051    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.152V 281.00ns 1.152V 301.00ns 1.050V 381.00ns 1.050V
Vi_052    i_052    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.195V 281.00ns 1.195V 301.00ns 1.050V 381.00ns 1.050V
Vi_053    i_053    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.258V 281.00ns 1.258V 301.00ns 1.050V 381.00ns 1.050V
Vi_054    i_054    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.188V 281.00ns 1.188V 301.00ns 1.050V 381.00ns 1.050V
Vi_055    i_055    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.228V 281.00ns 1.228V 301.00ns 1.050V 381.00ns 1.050V
Vi_056    i_056    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.313V 281.00ns 1.313V 301.00ns 1.050V 381.00ns 1.050V
Vi_057    i_057    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.087V 281.00ns 1.087V 301.00ns 1.050V 381.00ns 1.050V
Vi_058    i_058    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.146V 281.00ns 1.146V 301.00ns 1.050V 381.00ns 1.050V
Vi_059    i_059    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.166V 281.00ns 1.166V 301.00ns 1.050V 381.00ns 1.050V
Vi_060    i_060    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.199V 281.00ns 1.199V 301.00ns 1.050V 381.00ns 1.050V
Vi_061    i_061    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.274V 281.00ns 1.274V 301.00ns 1.050V 381.00ns 1.050V
Vi_062    i_062    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.200V 281.00ns 1.200V 301.00ns 1.050V 381.00ns 1.050V
Vi_063    i_063    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.208V 281.00ns 1.208V 301.00ns 1.050V 381.00ns 1.050V
Vi_064    i_064    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.350V 281.00ns 1.350V 301.00ns 1.050V 381.00ns 1.050V

* Vb_num: The bias voltage as pulse sequences

Vb_001    b_001    0    PWL 0.00ns 1.050V 1.00ns 1.050V 21.00ns 1.350V 281.00ns 1.350V 301.00ns 1.050V 381.00ns 1.050V
Vb_002    b_002    0    PWL 0.00ns 1.050V 11.00ns 1.050V 31.00ns 1.350V 291.00ns 1.350V 311.00ns 1.050V 391.00ns 1.050V
Vb_003    b_003    0    PWL 0.00ns 1.050V 21.00ns 1.050V 41.00ns 1.350V 301.00ns 1.350V 321.00ns 1.050V 401.00ns 1.050V

Ve        Ve       0    3
Vcc-      Vcc-     0    -5
Vcc+      Vcc+     0    5

* ============================ NN Parameters ==============================
* Parameters (weights and bias) naming convention: "Rl_i_j+" where:
*   R: Always "R" to inform Xyce it is a resistance
*   l: layer name, "h" for the hidden and output layers and "b" for the biases.
*   i: index of the weight of a neuron (start from 1)
*   j: index of the neuron (start from 1)
*   +: parameter polarity, + or -

* ----------------------------- Layers -----------------------------


* ----- Weights
* Layer 001

* Neuron 1
Rh001_001_001+    i_001    tia_h_in_001_001+    1210291.6352100708
Rh001_001_001-    i_001    tia_h_in_001_001-    51168.65281430691
Rh001_002_001+    i_002    tia_h_in_001_001+    1200681.639911038
Rh001_002_001-    i_002    tia_h_in_001_001-    42935.18402169747
Rh001_003_001+    i_003    tia_h_in_001_001+    111788.69723541531
Rh001_003_001-    i_003    tia_h_in_001_001-    1210338.5870977656
Rh001_004_001+    i_004    tia_h_in_001_001+    31464.77555878573
Rh001_004_001-    i_004    tia_h_in_001_001-    1189670.6792834178
Rh001_005_001+    i_005    tia_h_in_001_001+    26839.332857066107
Rh001_005_001-    i_005    tia_h_in_001_001-    1202835.956879755
Rh001_006_001+    i_006    tia_h_in_001_001+    33784.465329281455
Rh001_006_001-    i_006    tia_h_in_001_001-    1197439.4368922987
Rh001_007_001+    i_007    tia_h_in_001_001+    364953.3508063329
Rh001_007_001-    i_007    tia_h_in_001_001-    1201822.96121053
Rh001_008_001+    i_008    tia_h_in_001_001+    1192560.9752044221
Rh001_008_001-    i_008    tia_h_in_001_001-    306041.24189934117
Rh001_009_001+    i_009    tia_h_in_001_001+    224743.46620107105
Rh001_009_001-    i_009    tia_h_in_001_001-    1212004.6784558385
Rh001_010_001+    i_010    tia_h_in_001_001+    77198.6535396235
Rh001_010_001-    i_010    tia_h_in_001_001-    1211162.5447396631
Rh001_011_001+    i_011    tia_h_in_001_001+    36451.77495963238
Rh001_011_001-    i_011    tia_h_in_001_001-    1206367.1703335175
Rh001_012_001+    i_012    tia_h_in_001_001+    45350.7952886812
Rh001_012_001-    i_012    tia_h_in_001_001-    1199157.1564731402
Rh001_013_001+    i_013    tia_h_in_001_001+    67824.13848369135
Rh001_013_001-    i_013    tia_h_in_001_001-    1207495.533152037
Rh001_014_001+    i_014    tia_h_in_001_001+    1206173.407461235
Rh001_014_001-    i_014    tia_h_in_001_001-    362584.6976516861
Rh001_015_001+    i_015    tia_h_in_001_001+    1193226.6258906464
Rh001_015_001-    i_015    tia_h_in_001_001-    71231.64246786617
Rh001_016_001+    i_016    tia_h_in_001_001+    301733.13166284224
Rh001_016_001-    i_016    tia_h_in_001_001-    1210030.6710904636
Rh001_017_001+    i_017    tia_h_in_001_001+    1183783.2280535267
Rh001_017_001-    i_017    tia_h_in_001_001-    342090.1435229167
Rh001_018_001+    i_018    tia_h_in_001_001+    48377.55622527674
Rh001_018_001-    i_018    tia_h_in_001_001-    1190159.4465609612
Rh001_019_001+    i_019    tia_h_in_001_001+    64260.399002878956
Rh001_019_001-    i_019    tia_h_in_001_001-    1195975.075737011
Rh001_020_001+    i_020    tia_h_in_001_001+    31249.91296840082
Rh001_020_001-    i_020    tia_h_in_001_001-    1201078.946401058
Rh001_021_001+    i_021    tia_h_in_001_001+    103396.5141276146
Rh001_021_001-    i_021    tia_h_in_001_001-    1196156.702665817
Rh001_022_001+    i_022    tia_h_in_001_001+    1192938.8405307175
Rh001_022_001-    i_022    tia_h_in_001_001-    1024705.4573087909
Rh001_023_001+    i_023    tia_h_in_001_001+    596145.5392587036
Rh001_023_001-    i_023    tia_h_in_001_001-    1212107.30134822
Rh001_024_001+    i_024    tia_h_in_001_001+    1207513.5745084644
Rh001_024_001-    i_024    tia_h_in_001_001-    85686.2114856623
Rh001_025_001+    i_025    tia_h_in_001_001+    42474.13241256794
Rh001_025_001-    i_025    tia_h_in_001_001-    1190210.168892969
Rh001_026_001+    i_026    tia_h_in_001_001+    68010.08831596846
Rh001_026_001-    i_026    tia_h_in_001_001-    1186946.601905285
Rh001_027_001+    i_027    tia_h_in_001_001+    36064.10027850669
Rh001_027_001-    i_027    tia_h_in_001_001-    1189606.51384503
Rh001_028_001+    i_028    tia_h_in_001_001+    109148.44009011252
Rh001_028_001-    i_028    tia_h_in_001_001-    1217570.9400798022
Rh001_029_001+    i_029    tia_h_in_001_001+    1183178.407029879
Rh001_029_001-    i_029    tia_h_in_001_001-    130802.10507408819
Rh001_030_001+    i_030    tia_h_in_001_001+    1207810.0254754906
Rh001_030_001-    i_030    tia_h_in_001_001-    186176.91612118453
Rh001_031_001+    i_031    tia_h_in_001_001+    151705.1691848081
Rh001_031_001-    i_031    tia_h_in_001_001-    1202806.690945192
Rh001_032_001+    i_032    tia_h_in_001_001+    82199.72835941694
Rh001_032_001-    i_032    tia_h_in_001_001-    1182165.9987440365
Rh001_033_001+    i_033    tia_h_in_001_001+    85868.48089642792
Rh001_033_001-    i_033    tia_h_in_001_001-    1191037.1799881114
Rh001_034_001+    i_034    tia_h_in_001_001+    62548.89371967282
Rh001_034_001-    i_034    tia_h_in_001_001-    1184768.7889973202
Rh001_035_001+    i_035    tia_h_in_001_001+    147598.84571572972
Rh001_035_001-    i_035    tia_h_in_001_001-    1199932.7658445186
Rh001_036_001+    i_036    tia_h_in_001_001+    189440.55350674552
Rh001_036_001-    i_036    tia_h_in_001_001-    1175976.6591252568
Rh001_037_001+    i_037    tia_h_in_001_001+    262878.1350124112
Rh001_037_001-    i_037    tia_h_in_001_001-    1178978.5692287923
Rh001_038_001+    i_038    tia_h_in_001_001+    1208346.6672490975
Rh001_038_001-    i_038    tia_h_in_001_001-    354570.1171832381
Rh001_039_001+    i_039    tia_h_in_001_001+    745012.7576700136
Rh001_039_001-    i_039    tia_h_in_001_001-    1201564.2300286987
Rh001_040_001+    i_040    tia_h_in_001_001+    67226.74169754918
Rh001_040_001-    i_040    tia_h_in_001_001-    1187716.3829978292
Rh001_041_001+    i_041    tia_h_in_001_001+    56284.40770129444
Rh001_041_001-    i_041    tia_h_in_001_001-    1211825.20665206
Rh001_042_001+    i_042    tia_h_in_001_001+    1196915.1131744212
Rh001_042_001-    i_042    tia_h_in_001_001-    750503.7699444193
Rh001_043_001+    i_043    tia_h_in_001_001+    145652.96462084717
Rh001_043_001-    i_043    tia_h_in_001_001-    1194235.3647104267
Rh001_044_001+    i_044    tia_h_in_001_001+    1207554.4540835212
Rh001_044_001-    i_044    tia_h_in_001_001-    71015.11716845162
Rh001_045_001+    i_045    tia_h_in_001_001+    1189914.5381286195
Rh001_045_001-    i_045    tia_h_in_001_001-    1020311.7646466356
Rh001_046_001+    i_046    tia_h_in_001_001+    1199509.8030631982
Rh001_046_001-    i_046    tia_h_in_001_001-    398724.15352550993
Rh001_047_001+    i_047    tia_h_in_001_001+    77211.41890180997
Rh001_047_001-    i_047    tia_h_in_001_001-    1191862.3227856355
Rh001_048_001+    i_048    tia_h_in_001_001+    112037.05848665211
Rh001_048_001-    i_048    tia_h_in_001_001-    1199783.312552204
Rh001_049_001+    i_049    tia_h_in_001_001+    53106.60081790435
Rh001_049_001-    i_049    tia_h_in_001_001-    1181785.0518363973
Rh001_050_001+    i_050    tia_h_in_001_001+    51304.33328944812
Rh001_050_001-    i_050    tia_h_in_001_001-    1206887.708189354
Rh001_051_001+    i_051    tia_h_in_001_001+    212617.77102042915
Rh001_051_001-    i_051    tia_h_in_001_001-    1199923.9469474829
Rh001_052_001+    i_052    tia_h_in_001_001+    1194127.4813510953
Rh001_052_001-    i_052    tia_h_in_001_001-    404168.17792081647
Rh001_053_001+    i_053    tia_h_in_001_001+    1199177.596090793
Rh001_053_001-    i_053    tia_h_in_001_001-    147301.8972151937
Rh001_054_001+    i_054    tia_h_in_001_001+    1213637.2487882723
Rh001_054_001-    i_054    tia_h_in_001_001-    80932.47693338456
Rh001_055_001+    i_055    tia_h_in_001_001+    86606.5943969387
Rh001_055_001-    i_055    tia_h_in_001_001-    1197851.5995284826
Rh001_056_001+    i_056    tia_h_in_001_001+    1207248.7237827345
Rh001_056_001-    i_056    tia_h_in_001_001-    467332.8358282316
Rh001_057_001+    i_057    tia_h_in_001_001+    64338.07530044639
Rh001_057_001-    i_057    tia_h_in_001_001-    1191716.4052503044
Rh001_058_001+    i_058    tia_h_in_001_001+    218252.58902325408
Rh001_058_001-    i_058    tia_h_in_001_001-    1208439.6541885124
Rh001_059_001+    i_059    tia_h_in_001_001+    1205416.388758054
Rh001_059_001-    i_059    tia_h_in_001_001-    37043.46681150151
Rh001_060_001+    i_060    tia_h_in_001_001+    1197253.814517345
Rh001_060_001-    i_060    tia_h_in_001_001-    39157.48824973739
Rh001_061_001+    i_061    tia_h_in_001_001+    169464.05410001354
Rh001_061_001-    i_061    tia_h_in_001_001-    1210849.19115528
Rh001_062_001+    i_062    tia_h_in_001_001+    46872.15327338488
Rh001_062_001-    i_062    tia_h_in_001_001-    1209998.4715851697
Rh001_063_001+    i_063    tia_h_in_001_001+    32346.032277687947
Rh001_063_001-    i_063    tia_h_in_001_001-    1207274.230604788
Rh001_064_001+    i_064    tia_h_in_001_001+    37756.93972648275
Rh001_064_001-    i_064    tia_h_in_001_001-    1209293.7680338477

* Neuron 2
Rh001_001_002+    i_001    tia_h_in_001_002+    1200417.2208607257
Rh001_001_002-    i_001    tia_h_in_001_002-    69665.74350332802
Rh001_002_002+    i_002    tia_h_in_001_002+    1187356.5588811084
Rh001_002_002-    i_002    tia_h_in_001_002-    58513.70509059696
Rh001_003_002+    i_003    tia_h_in_001_002+    1197005.2622277378
Rh001_003_002-    i_003    tia_h_in_001_002-    369446.6924583857
Rh001_004_002+    i_004    tia_h_in_001_002+    1220884.3106261261
Rh001_004_002-    i_004    tia_h_in_001_002-    147809.2772272393
Rh001_005_002+    i_005    tia_h_in_001_002+    1017744.8347043344
Rh001_005_002-    i_005    tia_h_in_001_002-    1220297.1071118512
Rh001_006_002+    i_006    tia_h_in_001_002+    1178306.7010614849
Rh001_006_002-    i_006    tia_h_in_001_002-    76674.87761930327
Rh001_007_002+    i_007    tia_h_in_001_002+    1209313.3951743871
Rh001_007_002-    i_007    tia_h_in_001_002-    60944.14738191356
Rh001_008_002+    i_008    tia_h_in_001_002+    1215395.653411412
Rh001_008_002-    i_008    tia_h_in_001_002-    87633.11801305368
Rh001_009_002+    i_009    tia_h_in_001_002+    1206597.7217700975
Rh001_009_002-    i_009    tia_h_in_001_002-    48259.43474034904
Rh001_010_002+    i_010    tia_h_in_001_002+    49763.87031983808
Rh001_010_002-    i_010    tia_h_in_001_002-    1205777.3638753796
Rh001_011_002+    i_011    tia_h_in_001_002+    342768.09527480206
Rh001_011_002-    i_011    tia_h_in_001_002-    1213153.349808927
Rh001_012_002+    i_012    tia_h_in_001_002+    47692.753998457665
Rh001_012_002-    i_012    tia_h_in_001_002-    1201254.1991495655
Rh001_013_002+    i_013    tia_h_in_001_002+    112657.90540804053
Rh001_013_002-    i_013    tia_h_in_001_002-    1204518.2107751435
Rh001_014_002+    i_014    tia_h_in_001_002+    167863.68022435083
Rh001_014_002-    i_014    tia_h_in_001_002-    1191944.807823131
Rh001_015_002+    i_015    tia_h_in_001_002+    65642.50138018552
Rh001_015_002-    i_015    tia_h_in_001_002-    1195395.99314813
Rh001_016_002+    i_016    tia_h_in_001_002+    73064.0053424826
Rh001_016_002-    i_016    tia_h_in_001_002-    1205910.2034360308
Rh001_017_002+    i_017    tia_h_in_001_002+    35369.00624070411
Rh001_017_002-    i_017    tia_h_in_001_002-    1202478.4979455238
Rh001_018_002+    i_018    tia_h_in_001_002+    1193543.4471887057
Rh001_018_002-    i_018    tia_h_in_001_002-    1060208.895838077
Rh001_019_002+    i_019    tia_h_in_001_002+    127497.01239272056
Rh001_019_002-    i_019    tia_h_in_001_002-    1194643.5753544369
Rh001_020_002+    i_020    tia_h_in_001_002+    593376.7164217959
Rh001_020_002-    i_020    tia_h_in_001_002-    1200342.2209773164
Rh001_021_002+    i_021    tia_h_in_001_002+    101314.96750073957
Rh001_021_002-    i_021    tia_h_in_001_002-    1197392.7779992109
Rh001_022_002+    i_022    tia_h_in_001_002+    43769.26907270632
Rh001_022_002-    i_022    tia_h_in_001_002-    1193052.9867934731
Rh001_023_002+    i_023    tia_h_in_001_002+    32365.21254874418
Rh001_023_002-    i_023    tia_h_in_001_002-    1195338.4500740927
Rh001_024_002+    i_024    tia_h_in_001_002+    29957.651844513683
Rh001_024_002-    i_024    tia_h_in_001_002-    1194223.4606977617
Rh001_025_002+    i_025    tia_h_in_001_002+    61966.14310672303
Rh001_025_002-    i_025    tia_h_in_001_002-    1185549.6817385291
Rh001_026_002+    i_026    tia_h_in_001_002+    59373.32675029642
Rh001_026_002-    i_026    tia_h_in_001_002-    1224347.1283454194
Rh001_027_002+    i_027    tia_h_in_001_002+    1201745.42346362
Rh001_027_002-    i_027    tia_h_in_001_002-    490215.4491813436
Rh001_028_002+    i_028    tia_h_in_001_002+    1188027.2825148213
Rh001_028_002-    i_028    tia_h_in_001_002-    259724.1074431308
Rh001_029_002+    i_029    tia_h_in_001_002+    43273.43249891831
Rh001_029_002-    i_029    tia_h_in_001_002-    1201444.5734083373
Rh001_030_002+    i_030    tia_h_in_001_002+    90457.46088071147
Rh001_030_002-    i_030    tia_h_in_001_002-    1201968.1200838403
Rh001_031_002+    i_031    tia_h_in_001_002+    99392.72096167438
Rh001_031_002-    i_031    tia_h_in_001_002-    1203016.1364521256
Rh001_032_002+    i_032    tia_h_in_001_002+    135043.5503804024
Rh001_032_002-    i_032    tia_h_in_001_002-    1175960.8690476383
Rh001_033_002+    i_033    tia_h_in_001_002+    71835.33198855944
Rh001_033_002-    i_033    tia_h_in_001_002-    1206625.8540113957
Rh001_034_002+    i_034    tia_h_in_001_002+    63554.508790118234
Rh001_034_002-    i_034    tia_h_in_001_002-    1194275.7672627014
Rh001_035_002+    i_035    tia_h_in_001_002+    107172.49321766598
Rh001_035_002-    i_035    tia_h_in_001_002-    1201821.8356661848
Rh001_036_002+    i_036    tia_h_in_001_002+    260788.54313601248
Rh001_036_002-    i_036    tia_h_in_001_002-    1185370.5574523748
Rh001_037_002+    i_037    tia_h_in_001_002+    109761.30445877094
Rh001_037_002-    i_037    tia_h_in_001_002-    1189214.046414677
Rh001_038_002+    i_038    tia_h_in_001_002+    453279.47875770554
Rh001_038_002-    i_038    tia_h_in_001_002-    1213434.7366748035
Rh001_039_002+    i_039    tia_h_in_001_002+    1219560.6425165392
Rh001_039_002-    i_039    tia_h_in_001_002-    94010.5080593205
Rh001_040_002+    i_040    tia_h_in_001_002+    1210310.398449774
Rh001_040_002-    i_040    tia_h_in_001_002-    338782.0414377052
Rh001_041_002+    i_041    tia_h_in_001_002+    118012.8947159614
Rh001_041_002-    i_041    tia_h_in_001_002-    1192303.6223777398
Rh001_042_002+    i_042    tia_h_in_001_002+    68017.31122195367
Rh001_042_002-    i_042    tia_h_in_001_002-    1203688.4313094744
Rh001_043_002+    i_043    tia_h_in_001_002+    38920.35458624248
Rh001_043_002-    i_043    tia_h_in_001_002-    1204313.6498455354
Rh001_044_002+    i_044    tia_h_in_001_002+    63417.21444046644
Rh001_044_002-    i_044    tia_h_in_001_002-    1203946.279426887
Rh001_045_002+    i_045    tia_h_in_001_002+    1195239.5429126006
Rh001_045_002-    i_045    tia_h_in_001_002-    121793.25294028445
Rh001_046_002+    i_046    tia_h_in_001_002+    1223934.2463613376
Rh001_046_002-    i_046    tia_h_in_001_002-    100539.69549003265
Rh001_047_002+    i_047    tia_h_in_001_002+    439241.8365332938
Rh001_047_002-    i_047    tia_h_in_001_002-    1189499.789949707
Rh001_048_002+    i_048    tia_h_in_001_002+    246842.32288579678
Rh001_048_002-    i_048    tia_h_in_001_002-    1213257.9798868343
Rh001_049_002+    i_049    tia_h_in_001_002+    1201765.6442865497
Rh001_049_002-    i_049    tia_h_in_001_002-    243454.11122235618
Rh001_050_002+    i_050    tia_h_in_001_002+    196815.32139523813
Rh001_050_002-    i_050    tia_h_in_001_002-    1184491.6171497582
Rh001_051_002+    i_051    tia_h_in_001_002+    262780.8433604103
Rh001_051_002-    i_051    tia_h_in_001_002-    1206800.154061051
Rh001_052_002+    i_052    tia_h_in_001_002+    194142.33831210222
Rh001_052_002-    i_052    tia_h_in_001_002-    1194089.9567812204
Rh001_053_002+    i_053    tia_h_in_001_002+    258934.05497093848
Rh001_053_002-    i_053    tia_h_in_001_002-    1197833.502390502
Rh001_054_002+    i_054    tia_h_in_001_002+    62681.57959044636
Rh001_054_002-    i_054    tia_h_in_001_002-    1202779.3577636036
Rh001_055_002+    i_055    tia_h_in_001_002+    1195848.7828560825
Rh001_055_002-    i_055    tia_h_in_001_002-    779784.2191450045
Rh001_056_002+    i_056    tia_h_in_001_002+    1206898.5107095442
Rh001_056_002-    i_056    tia_h_in_001_002-    96558.85152466626
Rh001_057_002+    i_057    tia_h_in_001_002+    175614.514933384
Rh001_057_002-    i_057    tia_h_in_001_002-    1196084.71367332
Rh001_058_002+    i_058    tia_h_in_001_002+    171743.4538753305
Rh001_058_002-    i_058    tia_h_in_001_002-    1194078.080203219
Rh001_059_002+    i_059    tia_h_in_001_002+    1207307.9809218028
Rh001_059_002-    i_059    tia_h_in_001_002-    454331.4890493611
Rh001_060_002+    i_060    tia_h_in_001_002+    152129.26634818572
Rh001_060_002-    i_060    tia_h_in_001_002-    1192956.0527931624
Rh001_061_002+    i_061    tia_h_in_001_002+    45587.05078908326
Rh001_061_002-    i_061    tia_h_in_001_002-    1192936.4471043444
Rh001_062_002+    i_062    tia_h_in_001_002+    83546.31174456836
Rh001_062_002-    i_062    tia_h_in_001_002-    1199702.7736167214
Rh001_063_002+    i_063    tia_h_in_001_002+    57421.96848684801
Rh001_063_002-    i_063    tia_h_in_001_002-    1207623.1704315445
Rh001_064_002+    i_064    tia_h_in_001_002+    1204295.0522306385
Rh001_064_002-    i_064    tia_h_in_001_002-    451161.10337781336

* Neuron 3
Rh001_001_003+    i_001    tia_h_in_001_003+    1209601.3649939173
Rh001_001_003-    i_001    tia_h_in_001_003-    327294.18860198173
Rh001_002_003+    i_002    tia_h_in_001_003+    1221054.1250262533
Rh001_002_003-    i_002    tia_h_in_001_003-    1197890.2438092583
Rh001_003_003+    i_003    tia_h_in_001_003+    32549.509991452403
Rh001_003_003-    i_003    tia_h_in_001_003-    1200603.0739658433
Rh001_004_003+    i_004    tia_h_in_001_003+    20751.210611478597
Rh001_004_003-    i_004    tia_h_in_001_003-    1219199.1858830338
Rh001_005_003+    i_005    tia_h_in_001_003+    41789.98826017354
Rh001_005_003-    i_005    tia_h_in_001_003-    1199615.3281168665
Rh001_006_003+    i_006    tia_h_in_001_003+    247431.06685167385
Rh001_006_003-    i_006    tia_h_in_001_003-    1195928.3493361853
Rh001_007_003+    i_007    tia_h_in_001_003+    1195308.240580604
Rh001_007_003-    i_007    tia_h_in_001_003-    146552.88164031235
Rh001_008_003+    i_008    tia_h_in_001_003+    1203836.8943378218
Rh001_008_003-    i_008    tia_h_in_001_003-    36548.32421452358
Rh001_009_003+    i_009    tia_h_in_001_003+    77144.77287248825
Rh001_009_003-    i_009    tia_h_in_001_003-    1188732.1372869117
Rh001_010_003+    i_010    tia_h_in_001_003+    56551.71645010715
Rh001_010_003-    i_010    tia_h_in_001_003-    1196448.489639496
Rh001_011_003+    i_011    tia_h_in_001_003+    46596.39180606596
Rh001_011_003-    i_011    tia_h_in_001_003-    1189854.5739661814
Rh001_012_003+    i_012    tia_h_in_001_003+    408826.6173197493
Rh001_012_003-    i_012    tia_h_in_001_003-    1202204.030515012
Rh001_013_003+    i_013    tia_h_in_001_003+    159820.44966916577
Rh001_013_003-    i_013    tia_h_in_001_003-    1194144.5216376374
Rh001_014_003+    i_014    tia_h_in_001_003+    1197792.6400485195
Rh001_014_003-    i_014    tia_h_in_001_003-    235385.85654462426
Rh001_015_003+    i_015    tia_h_in_001_003+    1202653.015676351
Rh001_015_003-    i_015    tia_h_in_001_003-    153481.71920266852
Rh001_016_003+    i_016    tia_h_in_001_003+    353635.9408685428
Rh001_016_003-    i_016    tia_h_in_001_003-    1201638.10515824
Rh001_017_003+    i_017    tia_h_in_001_003+    79055.30754897301
Rh001_017_003-    i_017    tia_h_in_001_003-    1208517.8227166492
Rh001_018_003+    i_018    tia_h_in_001_003+    70636.06844104007
Rh001_018_003-    i_018    tia_h_in_001_003-    1197829.7934587928
Rh001_019_003+    i_019    tia_h_in_001_003+    37942.5044598723
Rh001_019_003-    i_019    tia_h_in_001_003-    1209685.6578987865
Rh001_020_003+    i_020    tia_h_in_001_003+    85562.318983712
Rh001_020_003-    i_020    tia_h_in_001_003-    1195696.6059759853
Rh001_021_003+    i_021    tia_h_in_001_003+    131993.77423733418
Rh001_021_003-    i_021    tia_h_in_001_003-    1189123.3980903833
Rh001_022_003+    i_022    tia_h_in_001_003+    1193593.788222867
Rh001_022_003-    i_022    tia_h_in_001_003-    138457.25836579726
Rh001_023_003+    i_023    tia_h_in_001_003+    1193666.983536222
Rh001_023_003-    i_023    tia_h_in_001_003-    323479.3786255748
Rh001_024_003+    i_024    tia_h_in_001_003+    1203438.1415196941
Rh001_024_003-    i_024    tia_h_in_001_003-    356791.5665755779
Rh001_025_003+    i_025    tia_h_in_001_003+    45652.15271792689
Rh001_025_003-    i_025    tia_h_in_001_003-    1189463.3413190201
Rh001_026_003+    i_026    tia_h_in_001_003+    68024.26661788598
Rh001_026_003-    i_026    tia_h_in_001_003-    1187035.24367002
Rh001_027_003+    i_027    tia_h_in_001_003+    86073.46825490968
Rh001_027_003-    i_027    tia_h_in_001_003-    1205524.7760753345
Rh001_028_003+    i_028    tia_h_in_001_003+    1193603.815610782
Rh001_028_003-    i_028    tia_h_in_001_003-    127067.56597049709
Rh001_029_003+    i_029    tia_h_in_001_003+    395195.2561483558
Rh001_029_003-    i_029    tia_h_in_001_003-    1202805.4252939261
Rh001_030_003+    i_030    tia_h_in_001_003+    434833.55494394636
Rh001_030_003-    i_030    tia_h_in_001_003-    1212989.895746753
Rh001_031_003+    i_031    tia_h_in_001_003+    94301.32777997339
Rh001_031_003-    i_031    tia_h_in_001_003-    1195083.9197456923
Rh001_032_003+    i_032    tia_h_in_001_003+    81444.54991139479
Rh001_032_003-    i_032    tia_h_in_001_003-    1197516.1172228765
Rh001_033_003+    i_033    tia_h_in_001_003+    65300.7630339216
Rh001_033_003-    i_033    tia_h_in_001_003-    1185150.103467083
Rh001_034_003+    i_034    tia_h_in_001_003+    59475.25390264315
Rh001_034_003-    i_034    tia_h_in_001_003-    1205062.8640467594
Rh001_035_003+    i_035    tia_h_in_001_003+    1187537.243179792
Rh001_035_003-    i_035    tia_h_in_001_003-    137062.49413143937
Rh001_036_003+    i_036    tia_h_in_001_003+    1200352.591821554
Rh001_036_003-    i_036    tia_h_in_001_003-    1077352.9014017323
Rh001_037_003+    i_037    tia_h_in_001_003+    209447.13090579052
Rh001_037_003-    i_037    tia_h_in_001_003-    1200835.6744043482
Rh001_038_003+    i_038    tia_h_in_001_003+    1196798.460697619
Rh001_038_003-    i_038    tia_h_in_001_003-    363553.50028255756
Rh001_039_003+    i_039    tia_h_in_001_003+    107204.54152162126
Rh001_039_003-    i_039    tia_h_in_001_003-    1206399.021378859
Rh001_040_003+    i_040    tia_h_in_001_003+    38853.13411959617
Rh001_040_003-    i_040    tia_h_in_001_003-    1202214.16869628
Rh001_041_003+    i_041    tia_h_in_001_003+    91568.43244549741
Rh001_041_003-    i_041    tia_h_in_001_003-    1205773.5462419188
Rh001_042_003+    i_042    tia_h_in_001_003+    150474.8609212363
Rh001_042_003-    i_042    tia_h_in_001_003-    1219877.9274123155
Rh001_043_003+    i_043    tia_h_in_001_003+    1214667.624336854
Rh001_043_003-    i_043    tia_h_in_001_003-    176923.81930306827
Rh001_044_003+    i_044    tia_h_in_001_003+    343010.7715408923
Rh001_044_003-    i_044    tia_h_in_001_003-    1198373.6176982205
Rh001_045_003+    i_045    tia_h_in_001_003+    321416.20917927695
Rh001_045_003-    i_045    tia_h_in_001_003-    1202577.530560169
Rh001_046_003+    i_046    tia_h_in_001_003+    106098.95961186528
Rh001_046_003-    i_046    tia_h_in_001_003-    1209690.0855613276
Rh001_047_003+    i_047    tia_h_in_001_003+    35984.42678728478
Rh001_047_003-    i_047    tia_h_in_001_003-    1212888.627552424
Rh001_048_003+    i_048    tia_h_in_001_003+    38980.945896850775
Rh001_048_003-    i_048    tia_h_in_001_003-    1198373.979641469
Rh001_049_003+    i_049    tia_h_in_001_003+    89122.10931681162
Rh001_049_003-    i_049    tia_h_in_001_003-    1206922.7126870896
Rh001_050_003+    i_050    tia_h_in_001_003+    1198959.9204324135
Rh001_050_003-    i_050    tia_h_in_001_003-    582312.5773721457
Rh001_051_003+    i_051    tia_h_in_001_003+    197476.5314582924
Rh001_051_003-    i_051    tia_h_in_001_003-    1202469.8395288724
Rh001_052_003+    i_052    tia_h_in_001_003+    1205086.6409881688
Rh001_052_003-    i_052    tia_h_in_001_003-    515727.56267862365
Rh001_053_003+    i_053    tia_h_in_001_003+    1189421.6424164674
Rh001_053_003-    i_053    tia_h_in_001_003-    152814.97848566645
Rh001_054_003+    i_054    tia_h_in_001_003+    467124.8997659458
Rh001_054_003-    i_054    tia_h_in_001_003-    1189233.4144861905
Rh001_055_003+    i_055    tia_h_in_001_003+    45711.83726464494
Rh001_055_003-    i_055    tia_h_in_001_003-    1208450.6337933675
Rh001_056_003+    i_056    tia_h_in_001_003+    83017.27875732383
Rh001_056_003-    i_056    tia_h_in_001_003-    1197977.8594593478
Rh001_057_003+    i_057    tia_h_in_001_003+    1204358.66132025
Rh001_057_003-    i_057    tia_h_in_001_003-    86264.55114914976
Rh001_058_003+    i_058    tia_h_in_001_003+    1212369.954378356
Rh001_058_003-    i_058    tia_h_in_001_003-    193350.52519369565
Rh001_059_003+    i_059    tia_h_in_001_003+    1204286.3218765955
Rh001_059_003-    i_059    tia_h_in_001_003-    68592.14236240079
Rh001_060_003+    i_060    tia_h_in_001_003+    1201485.514732849
Rh001_060_003-    i_060    tia_h_in_001_003-    100175.69088213182
Rh001_061_003+    i_061    tia_h_in_001_003+    56376.767688614294
Rh001_061_003-    i_061    tia_h_in_001_003-    1185398.3127214818
Rh001_062_003+    i_062    tia_h_in_001_003+    22877.369886737844
Rh001_062_003-    i_062    tia_h_in_001_003-    1203318.7516238282
Rh001_063_003+    i_063    tia_h_in_001_003+    56574.112903030094
Rh001_063_003-    i_063    tia_h_in_001_003-    1207781.7701021505
Rh001_064_003+    i_064    tia_h_in_001_003+    78873.1149507301
Rh001_064_003-    i_064    tia_h_in_001_003-    1195486.4870822697

* Neuron 4
Rh001_001_004+    i_001    tia_h_in_001_004+    146199.47734732158
Rh001_001_004-    i_001    tia_h_in_001_004-    1223620.4958296062
Rh001_002_004+    i_002    tia_h_in_001_004+    163806.3948705355
Rh001_002_004-    i_002    tia_h_in_001_004-    1210143.0344643588
Rh001_003_004+    i_003    tia_h_in_001_004+    113002.47189804746
Rh001_003_004-    i_003    tia_h_in_001_004-    1202570.6030504142
Rh001_004_004+    i_004    tia_h_in_001_004+    108823.54174328348
Rh001_004_004-    i_004    tia_h_in_001_004-    1172746.8309692224
Rh001_005_004+    i_005    tia_h_in_001_004+    1205771.7634874862
Rh001_005_004-    i_005    tia_h_in_001_004-    318933.8498738619
Rh001_006_004+    i_006    tia_h_in_001_004+    301670.5954114606
Rh001_006_004-    i_006    tia_h_in_001_004-    1199282.306632837
Rh001_007_004+    i_007    tia_h_in_001_004+    70729.38017144265
Rh001_007_004-    i_007    tia_h_in_001_004-    1205970.9082951676
Rh001_008_004+    i_008    tia_h_in_001_004+    98642.15236939728
Rh001_008_004-    i_008    tia_h_in_001_004-    1206755.4793648145
Rh001_009_004+    i_009    tia_h_in_001_004+    160659.2312796761
Rh001_009_004-    i_009    tia_h_in_001_004-    1204289.5792142258
Rh001_010_004+    i_010    tia_h_in_001_004+    855608.1528258296
Rh001_010_004-    i_010    tia_h_in_001_004-    1204333.3384375796
Rh001_011_004+    i_011    tia_h_in_001_004+    866940.2158941708
Rh001_011_004-    i_011    tia_h_in_001_004-    1193794.472148835
Rh001_012_004+    i_012    tia_h_in_001_004+    1189374.735024077
Rh001_012_004-    i_012    tia_h_in_001_004-    338649.7808959102
Rh001_013_004+    i_013    tia_h_in_001_004+    263270.17046423216
Rh001_013_004-    i_013    tia_h_in_001_004-    1195307.0772474029
Rh001_014_004+    i_014    tia_h_in_001_004+    103532.22756920161
Rh001_014_004-    i_014    tia_h_in_001_004-    1183099.6839109187
Rh001_015_004+    i_015    tia_h_in_001_004+    80800.6081392246
Rh001_015_004-    i_015    tia_h_in_001_004-    1217255.5097398406
Rh001_016_004+    i_016    tia_h_in_001_004+    93122.62495649424
Rh001_016_004-    i_016    tia_h_in_001_004-    1216421.9295987636
Rh001_017_004+    i_017    tia_h_in_001_004+    1200406.472218371
Rh001_017_004-    i_017    tia_h_in_001_004-    333921.3852531566
Rh001_018_004+    i_018    tia_h_in_001_004+    780286.0406151413
Rh001_018_004-    i_018    tia_h_in_001_004-    1196891.7994532192
Rh001_019_004+    i_019    tia_h_in_001_004+    191489.4374620262
Rh001_019_004-    i_019    tia_h_in_001_004-    1192465.4321020513
Rh001_020_004+    i_020    tia_h_in_001_004+    64751.30602415295
Rh001_020_004-    i_020    tia_h_in_001_004-    1213171.1194340028
Rh001_021_004+    i_021    tia_h_in_001_004+    125543.17011472686
Rh001_021_004-    i_021    tia_h_in_001_004-    1202762.669020136
Rh001_022_004+    i_022    tia_h_in_001_004+    234284.30406008576
Rh001_022_004-    i_022    tia_h_in_001_004-    1216931.5770054434
Rh001_023_004+    i_023    tia_h_in_001_004+    96590.48008020534
Rh001_023_004-    i_023    tia_h_in_001_004-    1195548.6195109873
Rh001_024_004+    i_024    tia_h_in_001_004+    317527.1087740822
Rh001_024_004-    i_024    tia_h_in_001_004-    1206157.8282191928
Rh001_025_004+    i_025    tia_h_in_001_004+    1188232.1033349214
Rh001_025_004-    i_025    tia_h_in_001_004-    1153273.4681548092
Rh001_026_004+    i_026    tia_h_in_001_004+    75174.89167225019
Rh001_026_004-    i_026    tia_h_in_001_004-    1190641.6110861595
Rh001_027_004+    i_027    tia_h_in_001_004+    384902.94024468795
Rh001_027_004-    i_027    tia_h_in_001_004-    1210021.799664389
Rh001_028_004+    i_028    tia_h_in_001_004+    200502.35157006962
Rh001_028_004-    i_028    tia_h_in_001_004-    1165153.5821202428
Rh001_029_004+    i_029    tia_h_in_001_004+    1208351.9460803878
Rh001_029_004-    i_029    tia_h_in_001_004-    252933.80260932766
Rh001_030_004+    i_030    tia_h_in_001_004+    79528.440274923
Rh001_030_004-    i_030    tia_h_in_001_004-    1195713.8135004311
Rh001_031_004+    i_031    tia_h_in_001_004+    75661.3268709642
Rh001_031_004-    i_031    tia_h_in_001_004-    1194056.3551529185
Rh001_032_004+    i_032    tia_h_in_001_004+    101744.44800627639
Rh001_032_004-    i_032    tia_h_in_001_004-    1197229.5249937503
Rh001_033_004+    i_033    tia_h_in_001_004+    1197428.9207981913
Rh001_033_004-    i_033    tia_h_in_001_004-    768897.3166214228
Rh001_034_004+    i_034    tia_h_in_001_004+    1204043.5433725836
Rh001_034_004-    i_034    tia_h_in_001_004-    260215.44112594915
Rh001_035_004+    i_035    tia_h_in_001_004+    1192541.1165212751
Rh001_035_004-    i_035    tia_h_in_001_004-    446536.7828296523
Rh001_036_004+    i_036    tia_h_in_001_004+    74155.55527601198
Rh001_036_004-    i_036    tia_h_in_001_004-    1193654.3345641254
Rh001_037_004+    i_037    tia_h_in_001_004+    90990.67386852858
Rh001_037_004-    i_037    tia_h_in_001_004-    1190244.7691766035
Rh001_038_004+    i_038    tia_h_in_001_004+    69784.30781031286
Rh001_038_004-    i_038    tia_h_in_001_004-    1197391.8105023452
Rh001_039_004+    i_039    tia_h_in_001_004+    88098.9460602006
Rh001_039_004-    i_039    tia_h_in_001_004-    1195017.8477406988
Rh001_040_004+    i_040    tia_h_in_001_004+    114186.83280329494
Rh001_040_004-    i_040    tia_h_in_001_004-    1195687.8936732365
Rh001_041_004+    i_041    tia_h_in_001_004+    148225.01273818105
Rh001_041_004-    i_041    tia_h_in_001_004-    1209024.639216987
Rh001_042_004+    i_042    tia_h_in_001_004+    1208889.192177162
Rh001_042_004-    i_042    tia_h_in_001_004-    558485.5689478066
Rh001_043_004+    i_043    tia_h_in_001_004+    1206566.17063879
Rh001_043_004-    i_043    tia_h_in_001_004-    391149.2736576416
Rh001_044_004+    i_044    tia_h_in_001_004+    1206113.1294223878
Rh001_044_004-    i_044    tia_h_in_001_004-    305175.1285203397
Rh001_045_004+    i_045    tia_h_in_001_004+    95016.82832205914
Rh001_045_004-    i_045    tia_h_in_001_004-    1196421.694675452
Rh001_046_004+    i_046    tia_h_in_001_004+    440127.40630624583
Rh001_046_004-    i_046    tia_h_in_001_004-    1196885.462699457
Rh001_047_004+    i_047    tia_h_in_001_004+    203365.7229706903
Rh001_047_004-    i_047    tia_h_in_001_004-    1191774.1710709669
Rh001_048_004+    i_048    tia_h_in_001_004+    704326.7290009125
Rh001_048_004-    i_048    tia_h_in_001_004-    1176379.928452084
Rh001_049_004+    i_049    tia_h_in_001_004+    203652.2933728354
Rh001_049_004-    i_049    tia_h_in_001_004-    1196415.9226217342
Rh001_050_004+    i_050    tia_h_in_001_004+    1212168.063629466
Rh001_050_004-    i_050    tia_h_in_001_004-    814008.2262846702
Rh001_051_004+    i_051    tia_h_in_001_004+    1040544.3136840536
Rh001_051_004-    i_051    tia_h_in_001_004-    1207699.2325778953
Rh001_052_004+    i_052    tia_h_in_001_004+    99322.93274260241
Rh001_052_004-    i_052    tia_h_in_001_004-    1202642.4923599903
Rh001_053_004+    i_053    tia_h_in_001_004+    245376.5243418519
Rh001_053_004-    i_053    tia_h_in_001_004-    1180684.674103638
Rh001_054_004+    i_054    tia_h_in_001_004+    81460.29374844821
Rh001_054_004-    i_054    tia_h_in_001_004-    1205370.767290666
Rh001_055_004+    i_055    tia_h_in_001_004+    260170.2378692564
Rh001_055_004-    i_055    tia_h_in_001_004-    1192806.4808499385
Rh001_056_004+    i_056    tia_h_in_001_004+    1198522.3189746004
Rh001_056_004-    i_056    tia_h_in_001_004-    609659.3037102632
Rh001_057_004+    i_057    tia_h_in_001_004+    195334.3216497564
Rh001_057_004-    i_057    tia_h_in_001_004-    1184580.1052511386
Rh001_058_004+    i_058    tia_h_in_001_004+    408847.30637199676
Rh001_058_004-    i_058    tia_h_in_001_004-    1203579.412423289
Rh001_059_004+    i_059    tia_h_in_001_004+    241535.7239407708
Rh001_059_004-    i_059    tia_h_in_001_004-    1205513.141718554
Rh001_060_004+    i_060    tia_h_in_001_004+    1193080.3212948288
Rh001_060_004-    i_060    tia_h_in_001_004-    310933.8489234788
Rh001_061_004+    i_061    tia_h_in_001_004+    84275.2645556302
Rh001_061_004-    i_061    tia_h_in_001_004-    1200397.734569875
Rh001_062_004+    i_062    tia_h_in_001_004+    1214500.0342548522
Rh001_062_004-    i_062    tia_h_in_001_004-    879749.8957371232
Rh001_063_004+    i_063    tia_h_in_001_004+    88055.53116080596
Rh001_063_004-    i_063    tia_h_in_001_004-    1200069.4294740115
Rh001_064_004+    i_064    tia_h_in_001_004+    94648.99411781685
Rh001_064_004-    i_064    tia_h_in_001_004-    1184870.6079859487

* Neuron 5
Rh001_001_005+    i_001    tia_h_in_001_005+    1202560.723755408
Rh001_001_005-    i_001    tia_h_in_001_005-    43707.1828466009
Rh001_002_005+    i_002    tia_h_in_001_005+    1208684.3143363749
Rh001_002_005-    i_002    tia_h_in_001_005-    39327.931531779985
Rh001_003_005+    i_003    tia_h_in_001_005+    1212498.3185762996
Rh001_003_005-    i_003    tia_h_in_001_005-    405989.1317022547
Rh001_004_005+    i_004    tia_h_in_001_005+    1188274.7051101155
Rh001_004_005-    i_004    tia_h_in_001_005-    128337.96547350436
Rh001_005_005+    i_005    tia_h_in_001_005+    1211651.2177614623
Rh001_005_005-    i_005    tia_h_in_001_005-    124426.4039399035
Rh001_006_005+    i_006    tia_h_in_001_005+    126861.43362597354
Rh001_006_005-    i_006    tia_h_in_001_005-    1192938.0714277276
Rh001_007_005+    i_007    tia_h_in_001_005+    1207972.2139065934
Rh001_007_005-    i_007    tia_h_in_001_005-    162054.59289835824
Rh001_008_005+    i_008    tia_h_in_001_005+    241709.90013821865
Rh001_008_005-    i_008    tia_h_in_001_005-    1181432.9482418601
Rh001_009_005+    i_009    tia_h_in_001_005+    107195.74222135493
Rh001_009_005-    i_009    tia_h_in_001_005-    1193539.003652277
Rh001_010_005+    i_010    tia_h_in_001_005+    26848.930653234456
Rh001_010_005-    i_010    tia_h_in_001_005-    1191141.7629344992
Rh001_011_005+    i_011    tia_h_in_001_005+    47817.53251423598
Rh001_011_005-    i_011    tia_h_in_001_005-    1189266.386972098
Rh001_012_005+    i_012    tia_h_in_001_005+    101549.91857463557
Rh001_012_005-    i_012    tia_h_in_001_005-    1200799.1830854614
Rh001_013_005+    i_013    tia_h_in_001_005+    65866.89417843019
Rh001_013_005-    i_013    tia_h_in_001_005-    1183478.2331361677
Rh001_014_005+    i_014    tia_h_in_001_005+    42087.90665034987
Rh001_014_005-    i_014    tia_h_in_001_005-    1200662.7379415308
Rh001_015_005+    i_015    tia_h_in_001_005+    42976.622690302866
Rh001_015_005-    i_015    tia_h_in_001_005-    1201846.3395171887
Rh001_016_005+    i_016    tia_h_in_001_005+    48737.77201655764
Rh001_016_005-    i_016    tia_h_in_001_005-    1195447.7951539746
Rh001_017_005+    i_017    tia_h_in_001_005+    227099.08712282465
Rh001_017_005-    i_017    tia_h_in_001_005-    1190213.8740925542
Rh001_018_005+    i_018    tia_h_in_001_005+    386247.40631990146
Rh001_018_005-    i_018    tia_h_in_001_005-    1190784.0694806247
Rh001_019_005+    i_019    tia_h_in_001_005+    48883.540938964
Rh001_019_005-    i_019    tia_h_in_001_005-    1187611.40969709
Rh001_020_005+    i_020    tia_h_in_001_005+    133372.06642723427
Rh001_020_005-    i_020    tia_h_in_001_005-    1203320.4120313644
Rh001_021_005+    i_021    tia_h_in_001_005+    535713.4465567424
Rh001_021_005-    i_021    tia_h_in_001_005-    1200730.0623211171
Rh001_022_005+    i_022    tia_h_in_001_005+    1202858.8584400974
Rh001_022_005-    i_022    tia_h_in_001_005-    112622.64968108204
Rh001_023_005+    i_023    tia_h_in_001_005+    1201809.9730788807
Rh001_023_005-    i_023    tia_h_in_001_005-    146131.42856929937
Rh001_024_005+    i_024    tia_h_in_001_005+    87116.52816160714
Rh001_024_005-    i_024    tia_h_in_001_005-    1195218.0830013303
Rh001_025_005+    i_025    tia_h_in_001_005+    133052.17594564846
Rh001_025_005-    i_025    tia_h_in_001_005-    1213805.959586019
Rh001_026_005+    i_026    tia_h_in_001_005+    82725.85397285181
Rh001_026_005-    i_026    tia_h_in_001_005-    1196825.106350579
Rh001_027_005+    i_027    tia_h_in_001_005+    83687.26510556866
Rh001_027_005-    i_027    tia_h_in_001_005-    1202021.4495554822
Rh001_028_005+    i_028    tia_h_in_001_005+    70182.44116045762
Rh001_028_005-    i_028    tia_h_in_001_005-    1187971.9130491314
Rh001_029_005+    i_029    tia_h_in_001_005+    197824.66109434678
Rh001_029_005-    i_029    tia_h_in_001_005-    1201564.5538953405
Rh001_030_005+    i_030    tia_h_in_001_005+    1206983.1367817533
Rh001_030_005-    i_030    tia_h_in_001_005-    231753.5243692904
Rh001_031_005+    i_031    tia_h_in_001_005+    76134.37991639276
Rh001_031_005-    i_031    tia_h_in_001_005-    1192389.7687033128
Rh001_032_005+    i_032    tia_h_in_001_005+    66892.84893816094
Rh001_032_005-    i_032    tia_h_in_001_005-    1209701.5415834303
Rh001_033_005+    i_033    tia_h_in_001_005+    1209907.5693282753
Rh001_033_005-    i_033    tia_h_in_001_005-    1119175.6379732804
Rh001_034_005+    i_034    tia_h_in_001_005+    1191007.845491469
Rh001_034_005-    i_034    tia_h_in_001_005-    121978.23864098622
Rh001_035_005+    i_035    tia_h_in_001_005+    447132.11376797216
Rh001_035_005-    i_035    tia_h_in_001_005-    1202034.1936147758
Rh001_036_005+    i_036    tia_h_in_001_005+    124441.80322829814
Rh001_036_005-    i_036    tia_h_in_001_005-    1204437.2499435325
Rh001_037_005+    i_037    tia_h_in_001_005+    128516.7185857361
Rh001_037_005-    i_037    tia_h_in_001_005-    1209929.5067307504
Rh001_038_005+    i_038    tia_h_in_001_005+    277417.3023002842
Rh001_038_005-    i_038    tia_h_in_001_005-    1203481.48730377
Rh001_039_005+    i_039    tia_h_in_001_005+    1211302.7684103276
Rh001_039_005-    i_039    tia_h_in_001_005-    705644.2181437536
Rh001_040_005+    i_040    tia_h_in_001_005+    89857.82311957907
Rh001_040_005-    i_040    tia_h_in_001_005-    1203302.975200914
Rh001_041_005+    i_041    tia_h_in_001_005+    91680.97825323013
Rh001_041_005-    i_041    tia_h_in_001_005-    1209123.7551198495
Rh001_042_005+    i_042    tia_h_in_001_005+    263457.47475665796
Rh001_042_005-    i_042    tia_h_in_001_005-    1199199.3497789933
Rh001_043_005+    i_043    tia_h_in_001_005+    1213040.2983640858
Rh001_043_005-    i_043    tia_h_in_001_005-    54616.6340235758
Rh001_044_005+    i_044    tia_h_in_001_005+    61185.34597431449
Rh001_044_005-    i_044    tia_h_in_001_005-    1205005.3613418692
Rh001_045_005+    i_045    tia_h_in_001_005+    50676.88171142378
Rh001_045_005-    i_045    tia_h_in_001_005-    1204835.1979621707
Rh001_046_005+    i_046    tia_h_in_001_005+    208435.96203910792
Rh001_046_005-    i_046    tia_h_in_001_005-    1199704.289875541
Rh001_047_005+    i_047    tia_h_in_001_005+    1206376.4928623317
Rh001_047_005-    i_047    tia_h_in_001_005-    58409.06778200628
Rh001_048_005+    i_048    tia_h_in_001_005+    1203461.8610085153
Rh001_048_005-    i_048    tia_h_in_001_005-    213411.6999411904
Rh001_049_005+    i_049    tia_h_in_001_005+    174462.27097273993
Rh001_049_005-    i_049    tia_h_in_001_005-    1210162.8859426011
Rh001_050_005+    i_050    tia_h_in_001_005+    112799.11649682271
Rh001_050_005-    i_050    tia_h_in_001_005-    1206262.0105123536
Rh001_051_005+    i_051    tia_h_in_001_005+    69653.1680453376
Rh001_051_005-    i_051    tia_h_in_001_005-    1191423.1688007247
Rh001_052_005+    i_052    tia_h_in_001_005+    1203104.0141406038
Rh001_052_005-    i_052    tia_h_in_001_005-    183867.90125342057
Rh001_053_005+    i_053    tia_h_in_001_005+    108096.62789225689
Rh001_053_005-    i_053    tia_h_in_001_005-    1192264.3212509349
Rh001_054_005+    i_054    tia_h_in_001_005+    48430.03101092702
Rh001_054_005-    i_054    tia_h_in_001_005-    1206222.3353668638
Rh001_055_005+    i_055    tia_h_in_001_005+    43696.01627999892
Rh001_055_005-    i_055    tia_h_in_001_005-    1201714.0327960008
Rh001_056_005+    i_056    tia_h_in_001_005+    1186613.6335099372
Rh001_056_005-    i_056    tia_h_in_001_005-    334325.7383209105
Rh001_057_005+    i_057    tia_h_in_001_005+    68876.96229254006
Rh001_057_005-    i_057    tia_h_in_001_005-    1204423.5480788846
Rh001_058_005+    i_058    tia_h_in_001_005+    49191.66617821317
Rh001_058_005-    i_058    tia_h_in_001_005-    1215598.4031608903
Rh001_059_005+    i_059    tia_h_in_001_005+    75627.7028478143
Rh001_059_005-    i_059    tia_h_in_001_005-    1187108.8688606245
Rh001_060_005+    i_060    tia_h_in_001_005+    118215.32273919528
Rh001_060_005-    i_060    tia_h_in_001_005-    1207799.783289332
Rh001_061_005+    i_061    tia_h_in_001_005+    1202243.5460059273
Rh001_061_005-    i_061    tia_h_in_001_005-    653954.4593995016
Rh001_062_005+    i_062    tia_h_in_001_005+    76862.7112711735
Rh001_062_005-    i_062    tia_h_in_001_005-    1199768.3655952788
Rh001_063_005+    i_063    tia_h_in_001_005+    32395.108224284322
Rh001_063_005-    i_063    tia_h_in_001_005-    1192585.9065701237
Rh001_064_005+    i_064    tia_h_in_001_005+    1218572.4316081065
Rh001_064_005-    i_064    tia_h_in_001_005-    78730.47828410321

* Neuron 6
Rh001_001_006+    i_001    tia_h_in_001_006+    845864.6308764452
Rh001_001_006-    i_001    tia_h_in_001_006-    1216998.1087114615
Rh001_002_006+    i_002    tia_h_in_001_006+    1193107.1101295024
Rh001_002_006-    i_002    tia_h_in_001_006-    476433.4323522136
Rh001_003_006+    i_003    tia_h_in_001_006+    1178951.4963400424
Rh001_003_006-    i_003    tia_h_in_001_006-    939202.028823833
Rh001_004_006+    i_004    tia_h_in_001_006+    1198094.9836906225
Rh001_004_006-    i_004    tia_h_in_001_006-    261791.64300005432
Rh001_005_006+    i_005    tia_h_in_001_006+    1206763.4904867967
Rh001_005_006-    i_005    tia_h_in_001_006-    565624.558993751
Rh001_006_006+    i_006    tia_h_in_001_006+    219181.1964645574
Rh001_006_006-    i_006    tia_h_in_001_006-    1195127.7331674488
Rh001_007_006+    i_007    tia_h_in_001_006+    77405.1176663109
Rh001_007_006-    i_007    tia_h_in_001_006-    1206950.1893882407
Rh001_008_006+    i_008    tia_h_in_001_006+    118467.52013889654
Rh001_008_006-    i_008    tia_h_in_001_006-    1205531.9012477263
Rh001_009_006+    i_009    tia_h_in_001_006+    1195904.749670415
Rh001_009_006-    i_009    tia_h_in_001_006-    654199.3160135852
Rh001_010_006+    i_010    tia_h_in_001_006+    1210481.8975819969
Rh001_010_006-    i_010    tia_h_in_001_006-    498554.51872410293
Rh001_011_006+    i_011    tia_h_in_001_006+    88436.11128110954
Rh001_011_006-    i_011    tia_h_in_001_006-    1207355.2391555547
Rh001_012_006+    i_012    tia_h_in_001_006+    1210853.6781020905
Rh001_012_006-    i_012    tia_h_in_001_006-    716370.824553757
Rh001_013_006+    i_013    tia_h_in_001_006+    176300.262735894
Rh001_013_006-    i_013    tia_h_in_001_006-    1209082.746044113
Rh001_014_006+    i_014    tia_h_in_001_006+    87963.45980957519
Rh001_014_006-    i_014    tia_h_in_001_006-    1179727.0233836134
Rh001_015_006+    i_015    tia_h_in_001_006+    365702.31050813996
Rh001_015_006-    i_015    tia_h_in_001_006-    1208988.454219105
Rh001_016_006+    i_016    tia_h_in_001_006+    168397.87902946043
Rh001_016_006-    i_016    tia_h_in_001_006-    1197980.2144592772
Rh001_017_006+    i_017    tia_h_in_001_006+    164087.34745984382
Rh001_017_006-    i_017    tia_h_in_001_006-    1200048.0997423013
Rh001_018_006+    i_018    tia_h_in_001_006+    214622.59742556032
Rh001_018_006-    i_018    tia_h_in_001_006-    1191183.9364490942
Rh001_019_006+    i_019    tia_h_in_001_006+    443245.4312731319
Rh001_019_006-    i_019    tia_h_in_001_006-    1190784.9205294126
Rh001_020_006+    i_020    tia_h_in_001_006+    1213487.6913179911
Rh001_020_006-    i_020    tia_h_in_001_006-    343488.01221066626
Rh001_021_006+    i_021    tia_h_in_001_006+    1192894.7676850592
Rh001_021_006-    i_021    tia_h_in_001_006-    450439.1573989979
Rh001_022_006+    i_022    tia_h_in_001_006+    503653.6612944337
Rh001_022_006-    i_022    tia_h_in_001_006-    1212333.742086252
Rh001_023_006+    i_023    tia_h_in_001_006+    63787.55770350132
Rh001_023_006-    i_023    tia_h_in_001_006-    1200851.5876450494
Rh001_024_006+    i_024    tia_h_in_001_006+    384726.1471632447
Rh001_024_006-    i_024    tia_h_in_001_006-    1204170.2876721693
Rh001_025_006+    i_025    tia_h_in_001_006+    1194482.9048749416
Rh001_025_006-    i_025    tia_h_in_001_006-    1205107.4577752936
Rh001_026_006+    i_026    tia_h_in_001_006+    110650.22221808598
Rh001_026_006-    i_026    tia_h_in_001_006-    1209696.1638278558
Rh001_027_006+    i_027    tia_h_in_001_006+    105399.14204654902
Rh001_027_006-    i_027    tia_h_in_001_006-    1217779.1640130666
Rh001_028_006+    i_028    tia_h_in_001_006+    85045.95638782796
Rh001_028_006-    i_028    tia_h_in_001_006-    1214466.1180226007
Rh001_029_006+    i_029    tia_h_in_001_006+    74023.13521078766
Rh001_029_006-    i_029    tia_h_in_001_006-    1202171.3582878315
Rh001_030_006+    i_030    tia_h_in_001_006+    84720.94430028145
Rh001_030_006-    i_030    tia_h_in_001_006-    1199783.5521041134
Rh001_031_006+    i_031    tia_h_in_001_006+    1201326.2392390133
Rh001_031_006-    i_031    tia_h_in_001_006-    273907.4104140101
Rh001_032_006+    i_032    tia_h_in_001_006+    128974.23906132854
Rh001_032_006-    i_032    tia_h_in_001_006-    1203304.729329019
Rh001_033_006+    i_033    tia_h_in_001_006+    80771.62631775439
Rh001_033_006-    i_033    tia_h_in_001_006-    1199204.2540884777
Rh001_034_006+    i_034    tia_h_in_001_006+    166645.5266486034
Rh001_034_006-    i_034    tia_h_in_001_006-    1186739.4741342827
Rh001_035_006+    i_035    tia_h_in_001_006+    663167.850937837
Rh001_035_006-    i_035    tia_h_in_001_006-    1195250.3223472335
Rh001_036_006+    i_036    tia_h_in_001_006+    65236.539259087935
Rh001_036_006-    i_036    tia_h_in_001_006-    1199101.2924213859
Rh001_037_006+    i_037    tia_h_in_001_006+    306114.3762727162
Rh001_037_006-    i_037    tia_h_in_001_006-    1189308.522808742
Rh001_038_006+    i_038    tia_h_in_001_006+    596912.8310044929
Rh001_038_006-    i_038    tia_h_in_001_006-    1193796.6594468465
Rh001_039_006+    i_039    tia_h_in_001_006+    1191993.1076576028
Rh001_039_006-    i_039    tia_h_in_001_006-    345368.0125108914
Rh001_040_006+    i_040    tia_h_in_001_006+    136682.5162700172
Rh001_040_006-    i_040    tia_h_in_001_006-    1192746.9227713821
Rh001_041_006+    i_041    tia_h_in_001_006+    91795.41063842484
Rh001_041_006-    i_041    tia_h_in_001_006-    1212739.3777831194
Rh001_042_006+    i_042    tia_h_in_001_006+    113301.3694808712
Rh001_042_006-    i_042    tia_h_in_001_006-    1206894.2380894618
Rh001_043_006+    i_043    tia_h_in_001_006+    117593.68976051138
Rh001_043_006-    i_043    tia_h_in_001_006-    1190816.2861230588
Rh001_044_006+    i_044    tia_h_in_001_006+    1179515.5777147508
Rh001_044_006-    i_044    tia_h_in_001_006-    605100.649137062
Rh001_045_006+    i_045    tia_h_in_001_006+    1199891.023096708
Rh001_045_006-    i_045    tia_h_in_001_006-    307728.01394138526
Rh001_046_006+    i_046    tia_h_in_001_006+    143753.91723029033
Rh001_046_006-    i_046    tia_h_in_001_006-    1191680.1461059216
Rh001_047_006+    i_047    tia_h_in_001_006+    66536.62094113964
Rh001_047_006-    i_047    tia_h_in_001_006-    1204585.161133347
Rh001_048_006+    i_048    tia_h_in_001_006+    84094.6406376752
Rh001_048_006-    i_048    tia_h_in_001_006-    1215262.2448896444
Rh001_049_006+    i_049    tia_h_in_001_006+    617833.8743333968
Rh001_049_006-    i_049    tia_h_in_001_006-    1213781.9983212925
Rh001_050_006+    i_050    tia_h_in_001_006+    179415.77113345798
Rh001_050_006-    i_050    tia_h_in_001_006-    1216303.7064792064
Rh001_051_006+    i_051    tia_h_in_001_006+    1198859.0979071402
Rh001_051_006-    i_051    tia_h_in_001_006-    667610.9044434804
Rh001_052_006+    i_052    tia_h_in_001_006+    413748.7163314338
Rh001_052_006-    i_052    tia_h_in_001_006-    1204288.687426396
Rh001_053_006+    i_053    tia_h_in_001_006+    118327.61668643742
Rh001_053_006-    i_053    tia_h_in_001_006-    1192905.1551415727
Rh001_054_006+    i_054    tia_h_in_001_006+    84272.32405242398
Rh001_054_006-    i_054    tia_h_in_001_006-    1207134.1744088666
Rh001_055_006+    i_055    tia_h_in_001_006+    69616.7496481491
Rh001_055_006-    i_055    tia_h_in_001_006-    1214265.0331228036
Rh001_056_006+    i_056    tia_h_in_001_006+    1212865.0548519052
Rh001_056_006-    i_056    tia_h_in_001_006-    329940.3092540897
Rh001_057_006+    i_057    tia_h_in_001_006+    77140.36043082083
Rh001_057_006-    i_057    tia_h_in_001_006-    1212398.741008476
Rh001_058_006+    i_058    tia_h_in_001_006+    1216010.2756571316
Rh001_058_006-    i_058    tia_h_in_001_006-    843004.5875271703
Rh001_059_006+    i_059    tia_h_in_001_006+    98362.5558635831
Rh001_059_006-    i_059    tia_h_in_001_006-    1195411.0317783777
Rh001_060_006+    i_060    tia_h_in_001_006+    69427.7845241144
Rh001_060_006-    i_060    tia_h_in_001_006-    1194014.8030521725
Rh001_061_006+    i_061    tia_h_in_001_006+    144325.7651807654
Rh001_061_006-    i_061    tia_h_in_001_006-    1213685.977964288
Rh001_062_006+    i_062    tia_h_in_001_006+    66152.38223094094
Rh001_062_006-    i_062    tia_h_in_001_006-    1189951.6517407512
Rh001_063_006+    i_063    tia_h_in_001_006+    1200853.8242342467
Rh001_063_006-    i_063    tia_h_in_001_006-    410258.36300174677
Rh001_064_006+    i_064    tia_h_in_001_006+    288638.0346368328
Rh001_064_006-    i_064    tia_h_in_001_006-    1197509.3203041905

* Neuron 7
Rh001_001_007+    i_001    tia_h_in_001_007+    68758.87788607097
Rh001_001_007-    i_001    tia_h_in_001_007-    1193174.042508079
Rh001_002_007+    i_002    tia_h_in_001_007+    186507.45795516451
Rh001_002_007-    i_002    tia_h_in_001_007-    1196353.3797587198
Rh001_003_007+    i_003    tia_h_in_001_007+    308096.19424722024
Rh001_003_007-    i_003    tia_h_in_001_007-    1185093.9321251363
Rh001_004_007+    i_004    tia_h_in_001_007+    51512.34956284944
Rh001_004_007-    i_004    tia_h_in_001_007-    1206601.918522757
Rh001_005_007+    i_005    tia_h_in_001_007+    82042.4162510496
Rh001_005_007-    i_005    tia_h_in_001_007-    1201732.2743105846
Rh001_006_007+    i_006    tia_h_in_001_007+    96874.09041951162
Rh001_006_007-    i_006    tia_h_in_001_007-    1191825.6452298237
Rh001_007_007+    i_007    tia_h_in_001_007+    65231.39691292692
Rh001_007_007-    i_007    tia_h_in_001_007-    1215915.489137927
Rh001_008_007+    i_008    tia_h_in_001_007+    70374.43732848804
Rh001_008_007-    i_008    tia_h_in_001_007-    1204972.3870421574
Rh001_009_007+    i_009    tia_h_in_001_007+    1207701.3261562479
Rh001_009_007-    i_009    tia_h_in_001_007-    59504.37509617964
Rh001_010_007+    i_010    tia_h_in_001_007+    1199684.128125527
Rh001_010_007-    i_010    tia_h_in_001_007-    227778.22450966772
Rh001_011_007+    i_011    tia_h_in_001_007+    50569.52717797444
Rh001_011_007-    i_011    tia_h_in_001_007-    1195612.9299760002
Rh001_012_007+    i_012    tia_h_in_001_007+    65239.44775219043
Rh001_012_007-    i_012    tia_h_in_001_007-    1203989.2577769833
Rh001_013_007+    i_013    tia_h_in_001_007+    134011.45776676614
Rh001_013_007-    i_013    tia_h_in_001_007-    1198340.6448219544
Rh001_014_007+    i_014    tia_h_in_001_007+    49368.723961987605
Rh001_014_007-    i_014    tia_h_in_001_007-    1224812.4293533072
Rh001_015_007+    i_015    tia_h_in_001_007+    92166.23586674365
Rh001_015_007-    i_015    tia_h_in_001_007-    1204581.739765853
Rh001_016_007+    i_016    tia_h_in_001_007+    48574.85056236842
Rh001_016_007-    i_016    tia_h_in_001_007-    1212527.3409338302
Rh001_017_007+    i_017    tia_h_in_001_007+    1194812.2155956288
Rh001_017_007-    i_017    tia_h_in_001_007-    190887.08782116254
Rh001_018_007+    i_018    tia_h_in_001_007+    1177378.5863197397
Rh001_018_007-    i_018    tia_h_in_001_007-    311220.3991773212
Rh001_019_007+    i_019    tia_h_in_001_007+    1206517.4566332065
Rh001_019_007-    i_019    tia_h_in_001_007-    80902.64009856428
Rh001_020_007+    i_020    tia_h_in_001_007+    215209.50535480445
Rh001_020_007-    i_020    tia_h_in_001_007-    1206635.6284556242
Rh001_021_007+    i_021    tia_h_in_001_007+    669442.2196630803
Rh001_021_007-    i_021    tia_h_in_001_007-    1199685.141433243
Rh001_022_007+    i_022    tia_h_in_001_007+    1197532.1043649327
Rh001_022_007-    i_022    tia_h_in_001_007-    126170.97974577532
Rh001_023_007+    i_023    tia_h_in_001_007+    189079.32821618865
Rh001_023_007-    i_023    tia_h_in_001_007-    1200232.8863494606
Rh001_024_007+    i_024    tia_h_in_001_007+    115462.29085335879
Rh001_024_007-    i_024    tia_h_in_001_007-    1214715.7307398338
Rh001_025_007+    i_025    tia_h_in_001_007+    74987.4551929745
Rh001_025_007-    i_025    tia_h_in_001_007-    1192091.9810818392
Rh001_026_007+    i_026    tia_h_in_001_007+    43102.67179148467
Rh001_026_007-    i_026    tia_h_in_001_007-    1182304.385101381
Rh001_027_007+    i_027    tia_h_in_001_007+    111084.94429755639
Rh001_027_007-    i_027    tia_h_in_001_007-    1208295.2117891195
Rh001_028_007+    i_028    tia_h_in_001_007+    916815.476950469
Rh001_028_007-    i_028    tia_h_in_001_007-    1201514.2649806023
Rh001_029_007+    i_029    tia_h_in_001_007+    1211607.0683387064
Rh001_029_007-    i_029    tia_h_in_001_007-    268325.3000640472
Rh001_030_007+    i_030    tia_h_in_001_007+    163236.9317856717
Rh001_030_007-    i_030    tia_h_in_001_007-    1195041.7217695143
Rh001_031_007+    i_031    tia_h_in_001_007+    653911.5030982088
Rh001_031_007-    i_031    tia_h_in_001_007-    1198440.7123315479
Rh001_032_007+    i_032    tia_h_in_001_007+    255111.78872913503
Rh001_032_007-    i_032    tia_h_in_001_007-    1199556.4173366714
Rh001_033_007+    i_033    tia_h_in_001_007+    108409.19187550509
Rh001_033_007-    i_033    tia_h_in_001_007-    1181233.870519071
Rh001_034_007+    i_034    tia_h_in_001_007+    57081.255550716734
Rh001_034_007-    i_034    tia_h_in_001_007-    1203453.3942417968
Rh001_035_007+    i_035    tia_h_in_001_007+    1211257.8455346439
Rh001_035_007-    i_035    tia_h_in_001_007-    69548.20232933464
Rh001_036_007+    i_036    tia_h_in_001_007+    175253.36632851514
Rh001_036_007-    i_036    tia_h_in_001_007-    1196352.9213845055
Rh001_037_007+    i_037    tia_h_in_001_007+    73195.69800434764
Rh001_037_007-    i_037    tia_h_in_001_007-    1206004.234872744
Rh001_038_007+    i_038    tia_h_in_001_007+    1199417.115179128
Rh001_038_007-    i_038    tia_h_in_001_007-    192980.76857455436
Rh001_039_007+    i_039    tia_h_in_001_007+    71167.97091478764
Rh001_039_007-    i_039    tia_h_in_001_007-    1186656.6185294096
Rh001_040_007+    i_040    tia_h_in_001_007+    1198858.358301505
Rh001_040_007-    i_040    tia_h_in_001_007-    297729.2055758448
Rh001_041_007+    i_041    tia_h_in_001_007+    113214.78810153386
Rh001_041_007-    i_041    tia_h_in_001_007-    1188758.5122189648
Rh001_042_007+    i_042    tia_h_in_001_007+    66467.066627001
Rh001_042_007-    i_042    tia_h_in_001_007-    1201555.8174742332
Rh001_043_007+    i_043    tia_h_in_001_007+    206351.01653482078
Rh001_043_007-    i_043    tia_h_in_001_007-    1198682.8685072856
Rh001_044_007+    i_044    tia_h_in_001_007+    101502.06647108048
Rh001_044_007-    i_044    tia_h_in_001_007-    1202107.5915147075
Rh001_045_007+    i_045    tia_h_in_001_007+    1201272.5008108087
Rh001_045_007-    i_045    tia_h_in_001_007-    107269.72085927252
Rh001_046_007+    i_046    tia_h_in_001_007+    125060.60275376875
Rh001_046_007-    i_046    tia_h_in_001_007-    1186286.8527463318
Rh001_047_007+    i_047    tia_h_in_001_007+    55749.268761996595
Rh001_047_007-    i_047    tia_h_in_001_007-    1216555.6437971264
Rh001_048_007+    i_048    tia_h_in_001_007+    90332.68377063125
Rh001_048_007-    i_048    tia_h_in_001_007-    1203568.2225211875
Rh001_049_007+    i_049    tia_h_in_001_007+    94007.01849605414
Rh001_049_007-    i_049    tia_h_in_001_007-    1189127.7919050448
Rh001_050_007+    i_050    tia_h_in_001_007+    94812.59819536011
Rh001_050_007-    i_050    tia_h_in_001_007-    1200430.559153083
Rh001_051_007+    i_051    tia_h_in_001_007+    35202.03164174331
Rh001_051_007-    i_051    tia_h_in_001_007-    1200145.7593091552
Rh001_052_007+    i_052    tia_h_in_001_007+    58570.48834163974
Rh001_052_007-    i_052    tia_h_in_001_007-    1184402.4132311551
Rh001_053_007+    i_053    tia_h_in_001_007+    44445.58691622723
Rh001_053_007-    i_053    tia_h_in_001_007-    1200688.8365310584
Rh001_054_007+    i_054    tia_h_in_001_007+    27909.887951825716
Rh001_054_007-    i_054    tia_h_in_001_007-    1205099.3607562678
Rh001_055_007+    i_055    tia_h_in_001_007+    39519.148933886085
Rh001_055_007-    i_055    tia_h_in_001_007-    1200686.290520718
Rh001_056_007+    i_056    tia_h_in_001_007+    62692.043703532654
Rh001_056_007-    i_056    tia_h_in_001_007-    1216026.016262201
Rh001_057_007+    i_057    tia_h_in_001_007+    70886.87605600587
Rh001_057_007-    i_057    tia_h_in_001_007-    1201491.3647728914
Rh001_058_007+    i_058    tia_h_in_001_007+    417654.17668574705
Rh001_058_007-    i_058    tia_h_in_001_007-    1200358.742646423
Rh001_059_007+    i_059    tia_h_in_001_007+    1207158.9236004762
Rh001_059_007-    i_059    tia_h_in_001_007-    140058.69414335804
Rh001_060_007+    i_060    tia_h_in_001_007+    1201984.644162158
Rh001_060_007-    i_060    tia_h_in_001_007-    237373.39592216798
Rh001_061_007+    i_061    tia_h_in_001_007+    74150.98894138091
Rh001_061_007-    i_061    tia_h_in_001_007-    1203042.4728234338
Rh001_062_007+    i_062    tia_h_in_001_007+    1201898.5471435878
Rh001_062_007-    i_062    tia_h_in_001_007-    39434.171423073996
Rh001_063_007+    i_063    tia_h_in_001_007+    1188859.4312747514
Rh001_063_007-    i_063    tia_h_in_001_007-    27955.166888121847
Rh001_064_007+    i_064    tia_h_in_001_007+    1191905.5158534907
Rh001_064_007-    i_064    tia_h_in_001_007-    39432.14479782238

* Neuron 8
Rh001_001_008+    i_001    tia_h_in_001_008+    1201129.4964671666
Rh001_001_008-    i_001    tia_h_in_001_008-    112119.3910963643
Rh001_002_008+    i_002    tia_h_in_001_008+    52083.92046151531
Rh001_002_008-    i_002    tia_h_in_001_008-    1204652.734628488
Rh001_003_008+    i_003    tia_h_in_001_008+    1196427.0492315812
Rh001_003_008-    i_003    tia_h_in_001_008-    383581.0507508921
Rh001_004_008+    i_004    tia_h_in_001_008+    462655.25844560436
Rh001_004_008-    i_004    tia_h_in_001_008-    1195505.3486698412
Rh001_005_008+    i_005    tia_h_in_001_008+    122770.58775957597
Rh001_005_008-    i_005    tia_h_in_001_008-    1200227.1553010102
Rh001_006_008+    i_006    tia_h_in_001_008+    60452.0475297893
Rh001_006_008-    i_006    tia_h_in_001_008-    1195655.680232562
Rh001_007_008+    i_007    tia_h_in_001_008+    95899.91433580019
Rh001_007_008-    i_007    tia_h_in_001_008-    1202961.1430461043
Rh001_008_008+    i_008    tia_h_in_001_008+    36796.71217816032
Rh001_008_008-    i_008    tia_h_in_001_008-    1194577.3467879118
Rh001_009_008+    i_009    tia_h_in_001_008+    80712.96162149789
Rh001_009_008-    i_009    tia_h_in_001_008-    1201801.6815326295
Rh001_010_008+    i_010    tia_h_in_001_008+    97065.13119576017
Rh001_010_008-    i_010    tia_h_in_001_008-    1191789.9589842746
Rh001_011_008+    i_011    tia_h_in_001_008+    56198.38557224075
Rh001_011_008-    i_011    tia_h_in_001_008-    1193130.2860325153
Rh001_012_008+    i_012    tia_h_in_001_008+    1210150.2986566871
Rh001_012_008-    i_012    tia_h_in_001_008-    68223.24681291709
Rh001_013_008+    i_013    tia_h_in_001_008+    257155.09657578915
Rh001_013_008-    i_013    tia_h_in_001_008-    1210555.9619661104
Rh001_014_008+    i_014    tia_h_in_001_008+    1199901.6067038293
Rh001_014_008-    i_014    tia_h_in_001_008-    203502.0868912715
Rh001_015_008+    i_015    tia_h_in_001_008+    1219495.14188728
Rh001_015_008-    i_015    tia_h_in_001_008-    170225.2781315353
Rh001_016_008+    i_016    tia_h_in_001_008+    181768.49792031955
Rh001_016_008-    i_016    tia_h_in_001_008-    1210725.3409180413
Rh001_017_008+    i_017    tia_h_in_001_008+    37060.764210904264
Rh001_017_008-    i_017    tia_h_in_001_008-    1203648.6180754066
Rh001_018_008+    i_018    tia_h_in_001_008+    64273.89171084315
Rh001_018_008-    i_018    tia_h_in_001_008-    1207311.4465634394
Rh001_019_008+    i_019    tia_h_in_001_008+    37759.16144993265
Rh001_019_008-    i_019    tia_h_in_001_008-    1206424.0424399746
Rh001_020_008+    i_020    tia_h_in_001_008+    35942.546351485114
Rh001_020_008-    i_020    tia_h_in_001_008-    1190662.259059156
Rh001_021_008+    i_021    tia_h_in_001_008+    69250.7322363113
Rh001_021_008-    i_021    tia_h_in_001_008-    1196494.2146462742
Rh001_022_008+    i_022    tia_h_in_001_008+    1197213.71055626
Rh001_022_008-    i_022    tia_h_in_001_008-    207988.6843588153
Rh001_023_008+    i_023    tia_h_in_001_008+    106765.2703649878
Rh001_023_008-    i_023    tia_h_in_001_008-    1204436.8268075301
Rh001_024_008+    i_024    tia_h_in_001_008+    1201185.496535608
Rh001_024_008-    i_024    tia_h_in_001_008-    59017.580147219815
Rh001_025_008+    i_025    tia_h_in_001_008+    130551.47480117796
Rh001_025_008-    i_025    tia_h_in_001_008-    1193091.741735301
Rh001_026_008+    i_026    tia_h_in_001_008+    1184995.8659416744
Rh001_026_008-    i_026    tia_h_in_001_008-    473031.2927100263
Rh001_027_008+    i_027    tia_h_in_001_008+    91868.99900325916
Rh001_027_008-    i_027    tia_h_in_001_008-    1188873.7925270316
Rh001_028_008+    i_028    tia_h_in_001_008+    46157.143722071654
Rh001_028_008-    i_028    tia_h_in_001_008-    1197008.8469591527
Rh001_029_008+    i_029    tia_h_in_001_008+    212304.84077268073
Rh001_029_008-    i_029    tia_h_in_001_008-    1201941.6843449469
Rh001_030_008+    i_030    tia_h_in_001_008+    147818.30584488873
Rh001_030_008-    i_030    tia_h_in_001_008-    1206010.8217940405
Rh001_031_008+    i_031    tia_h_in_001_008+    1207209.4593045493
Rh001_031_008-    i_031    tia_h_in_001_008-    204310.11770120636
Rh001_032_008+    i_032    tia_h_in_001_008+    241281.72411321744
Rh001_032_008-    i_032    tia_h_in_001_008-    1194946.4094551615
Rh001_033_008+    i_033    tia_h_in_001_008+    1210367.9147956194
Rh001_033_008-    i_033    tia_h_in_001_008-    1016339.9805317961
Rh001_034_008+    i_034    tia_h_in_001_008+    78269.60781484918
Rh001_034_008-    i_034    tia_h_in_001_008-    1185886.062831596
Rh001_035_008+    i_035    tia_h_in_001_008+    105337.71515290928
Rh001_035_008-    i_035    tia_h_in_001_008-    1198372.6565707065
Rh001_036_008+    i_036    tia_h_in_001_008+    1206264.9979276713
Rh001_036_008-    i_036    tia_h_in_001_008-    88946.06176732635
Rh001_037_008+    i_037    tia_h_in_001_008+    62132.88424476321
Rh001_037_008-    i_037    tia_h_in_001_008-    1206712.4215331688
Rh001_038_008+    i_038    tia_h_in_001_008+    58326.1187977379
Rh001_038_008-    i_038    tia_h_in_001_008-    1205510.7763496395
Rh001_039_008+    i_039    tia_h_in_001_008+    149126.66640793663
Rh001_039_008-    i_039    tia_h_in_001_008-    1192587.8354070603
Rh001_040_008+    i_040    tia_h_in_001_008+    52792.66060025162
Rh001_040_008-    i_040    tia_h_in_001_008-    1177801.6149033532
Rh001_041_008+    i_041    tia_h_in_001_008+    1198962.2721128087
Rh001_041_008-    i_041    tia_h_in_001_008-    431439.7061673553
Rh001_042_008+    i_042    tia_h_in_001_008+    1196751.0166513317
Rh001_042_008-    i_042    tia_h_in_001_008-    73496.34404179572
Rh001_043_008+    i_043    tia_h_in_001_008+    1200680.6381110575
Rh001_043_008-    i_043    tia_h_in_001_008-    212032.71453210985
Rh001_044_008+    i_044    tia_h_in_001_008+    1201204.8815737453
Rh001_044_008-    i_044    tia_h_in_001_008-    163157.67655925287
Rh001_045_008+    i_045    tia_h_in_001_008+    96336.7360510393
Rh001_045_008-    i_045    tia_h_in_001_008-    1209765.9584020243
Rh001_046_008+    i_046    tia_h_in_001_008+    39609.76197681253
Rh001_046_008-    i_046    tia_h_in_001_008-    1203969.509097205
Rh001_047_008+    i_047    tia_h_in_001_008+    63753.9755806608
Rh001_047_008-    i_047    tia_h_in_001_008-    1193062.0919436994
Rh001_048_008+    i_048    tia_h_in_001_008+    27609.07511479292
Rh001_048_008-    i_048    tia_h_in_001_008-    1209625.7891192075
Rh001_049_008+    i_049    tia_h_in_001_008+    547400.2255996935
Rh001_049_008-    i_049    tia_h_in_001_008-    1200986.9886231392
Rh001_050_008+    i_050    tia_h_in_001_008+    85931.7541753446
Rh001_050_008-    i_050    tia_h_in_001_008-    1181331.7644893664
Rh001_051_008+    i_051    tia_h_in_001_008+    114933.82636085575
Rh001_051_008-    i_051    tia_h_in_001_008-    1196125.1976397426
Rh001_052_008+    i_052    tia_h_in_001_008+    54687.9295588269
Rh001_052_008-    i_052    tia_h_in_001_008-    1203521.0518446937
Rh001_053_008+    i_053    tia_h_in_001_008+    91593.40226806444
Rh001_053_008-    i_053    tia_h_in_001_008-    1202615.6025969323
Rh001_054_008+    i_054    tia_h_in_001_008+    37723.59387307444
Rh001_054_008-    i_054    tia_h_in_001_008-    1214491.2630586172
Rh001_055_008+    i_055    tia_h_in_001_008+    31979.898680269696
Rh001_055_008-    i_055    tia_h_in_001_008-    1185581.9160520907
Rh001_056_008+    i_056    tia_h_in_001_008+    78625.92520984384
Rh001_056_008-    i_056    tia_h_in_001_008-    1193382.0095530918
Rh001_057_008+    i_057    tia_h_in_001_008+    177041.59591538078
Rh001_057_008-    i_057    tia_h_in_001_008-    1203554.0335500308
Rh001_058_008+    i_058    tia_h_in_001_008+    312862.8944574256
Rh001_058_008-    i_058    tia_h_in_001_008-    1191793.8040181252
Rh001_059_008+    i_059    tia_h_in_001_008+    101143.8950051382
Rh001_059_008-    i_059    tia_h_in_001_008-    1207406.3162906182
Rh001_060_008+    i_060    tia_h_in_001_008+    1209694.5543834516
Rh001_060_008-    i_060    tia_h_in_001_008-    39370.40602321295
Rh001_061_008+    i_061    tia_h_in_001_008+    1209008.7872442876
Rh001_061_008-    i_061    tia_h_in_001_008-    91129.38120262956
Rh001_062_008+    i_062    tia_h_in_001_008+    1200174.8053703427
Rh001_062_008-    i_062    tia_h_in_001_008-    48607.36729759377
Rh001_063_008+    i_063    tia_h_in_001_008+    1187741.7241866067
Rh001_063_008-    i_063    tia_h_in_001_008-    23475.496123385987
Rh001_064_008+    i_064    tia_h_in_001_008+    1184295.9009254535
Rh001_064_008-    i_064    tia_h_in_001_008-    24706.129569329347

* Neuron 9
Rh001_001_009+    i_001    tia_h_in_001_009+    74285.06253428178
Rh001_001_009-    i_001    tia_h_in_001_009-    1205243.6728800454
Rh001_002_009+    i_002    tia_h_in_001_009+    1206689.1220354894
Rh001_002_009-    i_002    tia_h_in_001_009-    103119.15567685389
Rh001_003_009+    i_003    tia_h_in_001_009+    247928.83703741152
Rh001_003_009-    i_003    tia_h_in_001_009-    1215551.45242302
Rh001_004_009+    i_004    tia_h_in_001_009+    91421.74699268723
Rh001_004_009-    i_004    tia_h_in_001_009-    1195031.6891899751
Rh001_005_009+    i_005    tia_h_in_001_009+    118606.27514667287
Rh001_005_009-    i_005    tia_h_in_001_009-    1202346.0380109327
Rh001_006_009+    i_006    tia_h_in_001_009+    74597.58880684772
Rh001_006_009-    i_006    tia_h_in_001_009-    1220582.84877127
Rh001_007_009+    i_007    tia_h_in_001_009+    83468.97819922678
Rh001_007_009-    i_007    tia_h_in_001_009-    1176790.3837180792
Rh001_008_009+    i_008    tia_h_in_001_009+    60594.91113730407
Rh001_008_009-    i_008    tia_h_in_001_009-    1204201.7108198605
Rh001_009_009+    i_009    tia_h_in_001_009+    70068.97874633042
Rh001_009_009-    i_009    tia_h_in_001_009-    1201208.055838817
Rh001_010_009+    i_010    tia_h_in_001_009+    1198263.0664142638
Rh001_010_009-    i_010    tia_h_in_001_009-    718565.0067595836
Rh001_011_009+    i_011    tia_h_in_001_009+    103069.49580586297
Rh001_011_009-    i_011    tia_h_in_001_009-    1205342.4136157762
Rh001_012_009+    i_012    tia_h_in_001_009+    57716.181285867024
Rh001_012_009-    i_012    tia_h_in_001_009-    1207870.6745080403
Rh001_013_009+    i_013    tia_h_in_001_009+    1194449.6992599806
Rh001_013_009-    i_013    tia_h_in_001_009-    750819.7869836257
Rh001_014_009+    i_014    tia_h_in_001_009+    273530.37625379785
Rh001_014_009-    i_014    tia_h_in_001_009-    1197919.6087452113
Rh001_015_009+    i_015    tia_h_in_001_009+    647223.4727252834
Rh001_015_009-    i_015    tia_h_in_001_009-    1204028.9794411184
Rh001_016_009+    i_016    tia_h_in_001_009+    1204316.021059089
Rh001_016_009-    i_016    tia_h_in_001_009-    62782.64765344049
Rh001_017_009+    i_017    tia_h_in_001_009+    1194903.5981799304
Rh001_017_009-    i_017    tia_h_in_001_009-    54627.04047807791
Rh001_018_009+    i_018    tia_h_in_001_009+    33266.575457151506
Rh001_018_009-    i_018    tia_h_in_001_009-    1219957.4642895209
Rh001_019_009+    i_019    tia_h_in_001_009+    100973.87390246069
Rh001_019_009-    i_019    tia_h_in_001_009-    1194843.7545184055
Rh001_020_009+    i_020    tia_h_in_001_009+    222561.96442450187
Rh001_020_009-    i_020    tia_h_in_001_009-    1203217.3915007785
Rh001_021_009+    i_021    tia_h_in_001_009+    1215001.8723245014
Rh001_021_009-    i_021    tia_h_in_001_009-    232112.12296771575
Rh001_022_009+    i_022    tia_h_in_001_009+    687684.3762037358
Rh001_022_009-    i_022    tia_h_in_001_009-    1208229.4802901344
Rh001_023_009+    i_023    tia_h_in_001_009+    138202.68041513808
Rh001_023_009-    i_023    tia_h_in_001_009-    1197521.3791886016
Rh001_024_009+    i_024    tia_h_in_001_009+    61938.04839859425
Rh001_024_009-    i_024    tia_h_in_001_009-    1220795.8281777694
Rh001_025_009+    i_025    tia_h_in_001_009+    1195176.639681572
Rh001_025_009-    i_025    tia_h_in_001_009-    49488.92687655423
Rh001_026_009+    i_026    tia_h_in_001_009+    113040.2864366423
Rh001_026_009-    i_026    tia_h_in_001_009-    1191334.1542228754
Rh001_027_009+    i_027    tia_h_in_001_009+    212024.918598664
Rh001_027_009-    i_027    tia_h_in_001_009-    1192672.568043796
Rh001_028_009+    i_028    tia_h_in_001_009+    97157.6212014991
Rh001_028_009-    i_028    tia_h_in_001_009-    1196602.4070387224
Rh001_029_009+    i_029    tia_h_in_001_009+    86923.05437694113
Rh001_029_009-    i_029    tia_h_in_001_009-    1215083.2219766162
Rh001_030_009+    i_030    tia_h_in_001_009+    85768.2909877223
Rh001_030_009-    i_030    tia_h_in_001_009-    1202961.8528743607
Rh001_031_009+    i_031    tia_h_in_001_009+    61147.91506369832
Rh001_031_009-    i_031    tia_h_in_001_009-    1190374.4119118166
Rh001_032_009+    i_032    tia_h_in_001_009+    46455.951358735365
Rh001_032_009-    i_032    tia_h_in_001_009-    1193399.9824188293
Rh001_033_009+    i_033    tia_h_in_001_009+    44423.50811930235
Rh001_033_009-    i_033    tia_h_in_001_009-    1179553.939063137
Rh001_034_009+    i_034    tia_h_in_001_009+    73656.34891676731
Rh001_034_009-    i_034    tia_h_in_001_009-    1209901.7924274092
Rh001_035_009+    i_035    tia_h_in_001_009+    1073945.8192500803
Rh001_035_009-    i_035    tia_h_in_001_009-    1207321.0558900603
Rh001_036_009+    i_036    tia_h_in_001_009+    116432.89265568455
Rh001_036_009-    i_036    tia_h_in_001_009-    1187737.5526261933
Rh001_037_009+    i_037    tia_h_in_001_009+    159128.20293494774
Rh001_037_009-    i_037    tia_h_in_001_009-    1207980.0282462058
Rh001_038_009+    i_038    tia_h_in_001_009+    90114.32406327006
Rh001_038_009-    i_038    tia_h_in_001_009-    1184710.523445554
Rh001_039_009+    i_039    tia_h_in_001_009+    149783.52330454098
Rh001_039_009-    i_039    tia_h_in_001_009-    1205867.7174594903
Rh001_040_009+    i_040    tia_h_in_001_009+    57914.925808395725
Rh001_040_009-    i_040    tia_h_in_001_009-    1186002.7056271532
Rh001_041_009+    i_041    tia_h_in_001_009+    38476.65640892563
Rh001_041_009-    i_041    tia_h_in_001_009-    1173736.9629624493
Rh001_042_009+    i_042    tia_h_in_001_009+    91603.69484040087
Rh001_042_009-    i_042    tia_h_in_001_009-    1204753.479606245
Rh001_043_009+    i_043    tia_h_in_001_009+    92979.1666461858
Rh001_043_009-    i_043    tia_h_in_001_009-    1199949.6833240301
Rh001_044_009+    i_044    tia_h_in_001_009+    44106.89135853649
Rh001_044_009-    i_044    tia_h_in_001_009-    1184389.836987967
Rh001_045_009+    i_045    tia_h_in_001_009+    38069.90072733478
Rh001_045_009-    i_045    tia_h_in_001_009-    1207470.0027250852
Rh001_046_009+    i_046    tia_h_in_001_009+    88919.97508106956
Rh001_046_009-    i_046    tia_h_in_001_009-    1216242.4153433726
Rh001_047_009+    i_047    tia_h_in_001_009+    48059.55422140856
Rh001_047_009-    i_047    tia_h_in_001_009-    1185865.4877871813
Rh001_048_009+    i_048    tia_h_in_001_009+    28837.646113496958
Rh001_048_009-    i_048    tia_h_in_001_009-    1200327.9781901566
Rh001_049_009+    i_049    tia_h_in_001_009+    226045.96866527176
Rh001_049_009-    i_049    tia_h_in_001_009-    1210117.156424355
Rh001_050_009+    i_050    tia_h_in_001_009+    90345.21900565192
Rh001_050_009-    i_050    tia_h_in_001_009-    1189937.3461514723
Rh001_051_009+    i_051    tia_h_in_001_009+    1196908.6468603127
Rh001_051_009-    i_051    tia_h_in_001_009-    96593.74183006553
Rh001_052_009+    i_052    tia_h_in_001_009+    229965.43931261048
Rh001_052_009-    i_052    tia_h_in_001_009-    1206116.3619834103
Rh001_053_009+    i_053    tia_h_in_001_009+    1186026.7497365004
Rh001_053_009-    i_053    tia_h_in_001_009-    268630.4197558994
Rh001_054_009+    i_054    tia_h_in_001_009+    145576.10333685484
Rh001_054_009-    i_054    tia_h_in_001_009-    1215690.3394818346
Rh001_055_009+    i_055    tia_h_in_001_009+    58359.78466847401
Rh001_055_009-    i_055    tia_h_in_001_009-    1189287.3262458304
Rh001_056_009+    i_056    tia_h_in_001_009+    1204242.493397722
Rh001_056_009-    i_056    tia_h_in_001_009-    166349.94539179065
Rh001_057_009+    i_057    tia_h_in_001_009+    1200614.731128201
Rh001_057_009-    i_057    tia_h_in_001_009-    333891.00982828037
Rh001_058_009+    i_058    tia_h_in_001_009+    1208982.621425589
Rh001_058_009-    i_058    tia_h_in_001_009-    193582.09426511533
Rh001_059_009+    i_059    tia_h_in_001_009+    88069.01551578629
Rh001_059_009-    i_059    tia_h_in_001_009-    1207342.1989109998
Rh001_060_009+    i_060    tia_h_in_001_009+    1192882.86321747
Rh001_060_009-    i_060    tia_h_in_001_009-    192888.18224312036
Rh001_061_009+    i_061    tia_h_in_001_009+    1219664.5769392184
Rh001_061_009-    i_061    tia_h_in_001_009-    84028.05444194276
Rh001_062_009+    i_062    tia_h_in_001_009+    1204525.9656496057
Rh001_062_009-    i_062    tia_h_in_001_009-    296514.47227776184
Rh001_063_009+    i_063    tia_h_in_001_009+    1208215.0579540962
Rh001_063_009-    i_063    tia_h_in_001_009-    36912.38309428906
Rh001_064_009+    i_064    tia_h_in_001_009+    1224677.931224334
Rh001_064_009-    i_064    tia_h_in_001_009-    21764.7514323996

* Neuron 10
Rh001_001_010+    i_001    tia_h_in_001_010+    79899.9639435505
Rh001_001_010-    i_001    tia_h_in_001_010-    1197912.1218745832
Rh001_002_010+    i_002    tia_h_in_001_010+    1183605.7129885224
Rh001_002_010-    i_002    tia_h_in_001_010-    386955.64852358674
Rh001_003_010+    i_003    tia_h_in_001_010+    124497.98527291749
Rh001_003_010-    i_003    tia_h_in_001_010-    1196071.2198405822
Rh001_004_010+    i_004    tia_h_in_001_010+    67548.79705366374
Rh001_004_010-    i_004    tia_h_in_001_010-    1211002.617176269
Rh001_005_010+    i_005    tia_h_in_001_010+    118376.38046096874
Rh001_005_010-    i_005    tia_h_in_001_010-    1197058.0940971675
Rh001_006_010+    i_006    tia_h_in_001_010+    106892.80129473929
Rh001_006_010-    i_006    tia_h_in_001_010-    1198735.5316386358
Rh001_007_010+    i_007    tia_h_in_001_010+    533974.3653441197
Rh001_007_010-    i_007    tia_h_in_001_010-    1209809.3852018823
Rh001_008_010+    i_008    tia_h_in_001_010+    145264.45761042126
Rh001_008_010-    i_008    tia_h_in_001_010-    1205310.259294876
Rh001_009_010+    i_009    tia_h_in_001_010+    135497.85429379647
Rh001_009_010-    i_009    tia_h_in_001_010-    1194167.845980387
Rh001_010_010+    i_010    tia_h_in_001_010+    108006.97755716674
Rh001_010_010-    i_010    tia_h_in_001_010-    1195920.852869479
Rh001_011_010+    i_011    tia_h_in_001_010+    96659.55061698574
Rh001_011_010-    i_011    tia_h_in_001_010-    1209448.2354927638
Rh001_012_010+    i_012    tia_h_in_001_010+    67907.63668475559
Rh001_012_010-    i_012    tia_h_in_001_010-    1210253.139273433
Rh001_013_010+    i_013    tia_h_in_001_010+    1203463.68402287
Rh001_013_010-    i_013    tia_h_in_001_010-    683699.9498411757
Rh001_014_010+    i_014    tia_h_in_001_010+    139724.68383681777
Rh001_014_010-    i_014    tia_h_in_001_010-    1215646.3348998758
Rh001_015_010+    i_015    tia_h_in_001_010+    390157.7693841823
Rh001_015_010-    i_015    tia_h_in_001_010-    1209743.428037183
Rh001_016_010+    i_016    tia_h_in_001_010+    1198933.179432567
Rh001_016_010-    i_016    tia_h_in_001_010-    588052.2327810093
Rh001_017_010+    i_017    tia_h_in_001_010+    161032.92605033898
Rh001_017_010-    i_017    tia_h_in_001_010-    1184920.489290224
Rh001_018_010+    i_018    tia_h_in_001_010+    1188517.8279962076
Rh001_018_010-    i_018    tia_h_in_001_010-    381179.39341979654
Rh001_019_010+    i_019    tia_h_in_001_010+    77366.23391922923
Rh001_019_010-    i_019    tia_h_in_001_010-    1216050.571058014
Rh001_020_010+    i_020    tia_h_in_001_010+    124252.84122094765
Rh001_020_010-    i_020    tia_h_in_001_010-    1193284.7460177373
Rh001_021_010+    i_021    tia_h_in_001_010+    456746.03872950707
Rh001_021_010-    i_021    tia_h_in_001_010-    1195805.848061215
Rh001_022_010+    i_022    tia_h_in_001_010+    86566.8929395673
Rh001_022_010-    i_022    tia_h_in_001_010-    1189932.1005380966
Rh001_023_010+    i_023    tia_h_in_001_010+    1202061.456255685
Rh001_023_010-    i_023    tia_h_in_001_010-    307939.3642251136
Rh001_024_010+    i_024    tia_h_in_001_010+    281056.6642192513
Rh001_024_010-    i_024    tia_h_in_001_010-    1188198.1838460173
Rh001_025_010+    i_025    tia_h_in_001_010+    191833.26743188745
Rh001_025_010-    i_025    tia_h_in_001_010-    1197246.8173257343
Rh001_026_010+    i_026    tia_h_in_001_010+    1198090.6863603943
Rh001_026_010-    i_026    tia_h_in_001_010-    418792.9272823509
Rh001_027_010+    i_027    tia_h_in_001_010+    815818.7121254747
Rh001_027_010-    i_027    tia_h_in_001_010-    1196677.138709335
Rh001_028_010+    i_028    tia_h_in_001_010+    180786.52218373708
Rh001_028_010-    i_028    tia_h_in_001_010-    1200051.401345589
Rh001_029_010+    i_029    tia_h_in_001_010+    72244.24931255907
Rh001_029_010-    i_029    tia_h_in_001_010-    1208273.8843212642
Rh001_030_010+    i_030    tia_h_in_001_010+    63736.09183586277
Rh001_030_010-    i_030    tia_h_in_001_010-    1191429.8194016104
Rh001_031_010+    i_031    tia_h_in_001_010+    79525.80862524959
Rh001_031_010-    i_031    tia_h_in_001_010-    1189991.697753398
Rh001_032_010+    i_032    tia_h_in_001_010+    595349.0360349328
Rh001_032_010-    i_032    tia_h_in_001_010-    1190335.4506531183
Rh001_033_010+    i_033    tia_h_in_001_010+    980201.1519522761
Rh001_033_010-    i_033    tia_h_in_001_010-    1205418.7354649198
Rh001_034_010+    i_034    tia_h_in_001_010+    67321.72295535683
Rh001_034_010-    i_034    tia_h_in_001_010-    1196924.26068127
Rh001_035_010+    i_035    tia_h_in_001_010+    99186.30804078042
Rh001_035_010-    i_035    tia_h_in_001_010-    1190114.7174295345
Rh001_036_010+    i_036    tia_h_in_001_010+    139638.20271935518
Rh001_036_010-    i_036    tia_h_in_001_010-    1196564.3367903864
Rh001_037_010+    i_037    tia_h_in_001_010+    123728.96621858777
Rh001_037_010-    i_037    tia_h_in_001_010-    1210191.6847555893
Rh001_038_010+    i_038    tia_h_in_001_010+    1214173.5600476232
Rh001_038_010-    i_038    tia_h_in_001_010-    514984.8932031624
Rh001_039_010+    i_039    tia_h_in_001_010+    250937.10198677384
Rh001_039_010-    i_039    tia_h_in_001_010-    1193763.4307261535
Rh001_040_010+    i_040    tia_h_in_001_010+    64741.74869718933
Rh001_040_010-    i_040    tia_h_in_001_010-    1194871.715628593
Rh001_041_010+    i_041    tia_h_in_001_010+    211888.90730614547
Rh001_041_010-    i_041    tia_h_in_001_010-    1205896.7159570472
Rh001_042_010+    i_042    tia_h_in_001_010+    154337.1699259646
Rh001_042_010-    i_042    tia_h_in_001_010-    1207270.627092607
Rh001_043_010+    i_043    tia_h_in_001_010+    1182905.382431131
Rh001_043_010-    i_043    tia_h_in_001_010-    445873.3490120663
Rh001_044_010+    i_044    tia_h_in_001_010+    518108.42170039885
Rh001_044_010-    i_044    tia_h_in_001_010-    1200459.6050675514
Rh001_045_010+    i_045    tia_h_in_001_010+    148081.07447192768
Rh001_045_010-    i_045    tia_h_in_001_010-    1187121.9957948362
Rh001_046_010+    i_046    tia_h_in_001_010+    721856.2610373073
Rh001_046_010-    i_046    tia_h_in_001_010-    1200876.394720452
Rh001_047_010+    i_047    tia_h_in_001_010+    171496.5076997374
Rh001_047_010-    i_047    tia_h_in_001_010-    1214547.1350171966
Rh001_048_010+    i_048    tia_h_in_001_010+    92329.99220876372
Rh001_048_010-    i_048    tia_h_in_001_010-    1182292.6964765496
Rh001_049_010+    i_049    tia_h_in_001_010+    1195968.9149027616
Rh001_049_010-    i_049    tia_h_in_001_010-    298973.14758485893
Rh001_050_010+    i_050    tia_h_in_001_010+    104194.20841412326
Rh001_050_010-    i_050    tia_h_in_001_010-    1223135.181295817
Rh001_051_010+    i_051    tia_h_in_001_010+    875259.1278831896
Rh001_051_010-    i_051    tia_h_in_001_010-    1212931.2074580807
Rh001_052_010+    i_052    tia_h_in_001_010+    368225.34412185254
Rh001_052_010-    i_052    tia_h_in_001_010-    1176496.959284545
Rh001_053_010+    i_053    tia_h_in_001_010+    97625.36908762276
Rh001_053_010-    i_053    tia_h_in_001_010-    1206999.6870606919
Rh001_054_010+    i_054    tia_h_in_001_010+    70203.85902106001
Rh001_054_010-    i_054    tia_h_in_001_010-    1190607.9762457826
Rh001_055_010+    i_055    tia_h_in_001_010+    225705.68843016573
Rh001_055_010-    i_055    tia_h_in_001_010-    1211600.5666899602
Rh001_056_010+    i_056    tia_h_in_001_010+    309282.83971641207
Rh001_056_010-    i_056    tia_h_in_001_010-    1204432.1726506765
Rh001_057_010+    i_057    tia_h_in_001_010+    1187140.9120047716
Rh001_057_010-    i_057    tia_h_in_001_010-    343465.21057390654
Rh001_058_010+    i_058    tia_h_in_001_010+    440322.179720827
Rh001_058_010-    i_058    tia_h_in_001_010-    1197403.7006302276
Rh001_059_010+    i_059    tia_h_in_001_010+    1200094.4484732829
Rh001_059_010-    i_059    tia_h_in_001_010-    397936.4481101627
Rh001_060_010+    i_060    tia_h_in_001_010+    201478.4963987706
Rh001_060_010-    i_060    tia_h_in_001_010-    1212789.3980645856
Rh001_061_010+    i_061    tia_h_in_001_010+    113852.0597950538
Rh001_061_010-    i_061    tia_h_in_001_010-    1203581.0729055745
Rh001_062_010+    i_062    tia_h_in_001_010+    1180432.8790023401
Rh001_062_010-    i_062    tia_h_in_001_010-    322848.6143477508
Rh001_063_010+    i_063    tia_h_in_001_010+    68376.17272893347
Rh001_063_010-    i_063    tia_h_in_001_010-    1175388.5468010819
Rh001_064_010+    i_064    tia_h_in_001_010+    81372.78184416814
Rh001_064_010-    i_064    tia_h_in_001_010-    1216705.0225051832

* Neuron 11
Rh001_001_011+    i_001    tia_h_in_001_011+    1190285.5629896175
Rh001_001_011-    i_001    tia_h_in_001_011-    22286.98741348407
Rh001_002_011+    i_002    tia_h_in_001_011+    1212457.8369243585
Rh001_002_011-    i_002    tia_h_in_001_011-    53306.40196785678
Rh001_003_011+    i_003    tia_h_in_001_011+    1213259.7101826728
Rh001_003_011-    i_003    tia_h_in_001_011-    62850.74677943571
Rh001_004_011+    i_004    tia_h_in_001_011+    1190124.119979256
Rh001_004_011-    i_004    tia_h_in_001_011-    52703.327576446136
Rh001_005_011+    i_005    tia_h_in_001_011+    1205914.8532474004
Rh001_005_011-    i_005    tia_h_in_001_011-    87457.41363813453
Rh001_006_011+    i_006    tia_h_in_001_011+    1206046.6932927324
Rh001_006_011-    i_006    tia_h_in_001_011-    59932.194680337365
Rh001_007_011+    i_007    tia_h_in_001_011+    94117.31371157344
Rh001_007_011-    i_007    tia_h_in_001_011-    1186108.1438780404
Rh001_008_011+    i_008    tia_h_in_001_011+    153565.68012170258
Rh001_008_011-    i_008    tia_h_in_001_011-    1196312.6879024717
Rh001_009_011+    i_009    tia_h_in_001_011+    45416.09823065471
Rh001_009_011-    i_009    tia_h_in_001_011-    1196664.6581376905
Rh001_010_011+    i_010    tia_h_in_001_011+    47080.37930994127
Rh001_010_011-    i_010    tia_h_in_001_011-    1214071.33858334
Rh001_011_011+    i_011    tia_h_in_001_011+    35867.90669460493
Rh001_011_011-    i_011    tia_h_in_001_011-    1190948.7240564027
Rh001_012_011+    i_012    tia_h_in_001_011+    38489.21440962862
Rh001_012_011-    i_012    tia_h_in_001_011-    1201917.2328089003
Rh001_013_011+    i_013    tia_h_in_001_011+    84773.19538960126
Rh001_013_011-    i_013    tia_h_in_001_011-    1203419.0882387392
Rh001_014_011+    i_014    tia_h_in_001_011+    173926.27233324051
Rh001_014_011-    i_014    tia_h_in_001_011-    1208332.9658128878
Rh001_015_011+    i_015    tia_h_in_001_011+    1206064.6025449592
Rh001_015_011-    i_015    tia_h_in_001_011-    343203.8723961818
Rh001_016_011+    i_016    tia_h_in_001_011+    369887.7921164801
Rh001_016_011-    i_016    tia_h_in_001_011-    1210602.4568541
Rh001_017_011+    i_017    tia_h_in_001_011+    45450.34518685968
Rh001_017_011-    i_017    tia_h_in_001_011-    1219220.1179419416
Rh001_018_011+    i_018    tia_h_in_001_011+    42651.08251678185
Rh001_018_011-    i_018    tia_h_in_001_011-    1203383.6881985771
Rh001_019_011+    i_019    tia_h_in_001_011+    1205360.3738605788
Rh001_019_011-    i_019    tia_h_in_001_011-    481910.9281148014
Rh001_020_011+    i_020    tia_h_in_001_011+    51418.228313597916
Rh001_020_011-    i_020    tia_h_in_001_011-    1209623.5333974538
Rh001_021_011+    i_021    tia_h_in_001_011+    31210.696623937838
Rh001_021_011-    i_021    tia_h_in_001_011-    1194358.2124921302
Rh001_022_011+    i_022    tia_h_in_001_011+    85988.83826442309
Rh001_022_011-    i_022    tia_h_in_001_011-    1197602.916021246
Rh001_023_011+    i_023    tia_h_in_001_011+    139668.27421148855
Rh001_023_011-    i_023    tia_h_in_001_011-    1207383.3310248416
Rh001_024_011+    i_024    tia_h_in_001_011+    99782.0654479711
Rh001_024_011-    i_024    tia_h_in_001_011-    1192556.3109923238
Rh001_025_011+    i_025    tia_h_in_001_011+    60622.8110168638
Rh001_025_011-    i_025    tia_h_in_001_011-    1214617.830941347
Rh001_026_011+    i_026    tia_h_in_001_011+    1214726.319642008
Rh001_026_011-    i_026    tia_h_in_001_011-    153939.01503505986
Rh001_027_011+    i_027    tia_h_in_001_011+    151016.7042366815
Rh001_027_011-    i_027    tia_h_in_001_011-    1207504.7015968051
Rh001_028_011+    i_028    tia_h_in_001_011+    84224.92072377795
Rh001_028_011-    i_028    tia_h_in_001_011-    1199010.2555605415
Rh001_029_011+    i_029    tia_h_in_001_011+    98956.61190965757
Rh001_029_011-    i_029    tia_h_in_001_011-    1180775.5869041358
Rh001_030_011+    i_030    tia_h_in_001_011+    79199.99906290941
Rh001_030_011-    i_030    tia_h_in_001_011-    1194023.806603264
Rh001_031_011+    i_031    tia_h_in_001_011+    58164.507191532946
Rh001_031_011-    i_031    tia_h_in_001_011-    1200910.086190184
Rh001_032_011+    i_032    tia_h_in_001_011+    83118.30848185184
Rh001_032_011-    i_032    tia_h_in_001_011-    1198424.3203593832
Rh001_033_011+    i_033    tia_h_in_001_011+    183128.8282619926
Rh001_033_011-    i_033    tia_h_in_001_011-    1204793.5230185443
Rh001_034_011+    i_034    tia_h_in_001_011+    133542.336208494
Rh001_034_011-    i_034    tia_h_in_001_011-    1199848.4417488836
Rh001_035_011+    i_035    tia_h_in_001_011+    97939.51730824471
Rh001_035_011-    i_035    tia_h_in_001_011-    1206841.883721404
Rh001_036_011+    i_036    tia_h_in_001_011+    1215470.2439969413
Rh001_036_011-    i_036    tia_h_in_001_011-    71109.12517374782
Rh001_037_011+    i_037    tia_h_in_001_011+    163570.6281162357
Rh001_037_011-    i_037    tia_h_in_001_011-    1204780.5805981671
Rh001_038_011+    i_038    tia_h_in_001_011+    66551.13098676859
Rh001_038_011-    i_038    tia_h_in_001_011-    1199115.916247561
Rh001_039_011+    i_039    tia_h_in_001_011+    67552.88385516174
Rh001_039_011-    i_039    tia_h_in_001_011-    1199963.9160110722
Rh001_040_011+    i_040    tia_h_in_001_011+    1209433.3324919504
Rh001_040_011-    i_040    tia_h_in_001_011-    100620.86488869088
Rh001_041_011+    i_041    tia_h_in_001_011+    89826.59350213523
Rh001_041_011-    i_041    tia_h_in_001_011-    1212414.2366957308
Rh001_042_011+    i_042    tia_h_in_001_011+    136542.58684820827
Rh001_042_011-    i_042    tia_h_in_001_011-    1205051.4792553838
Rh001_043_011+    i_043    tia_h_in_001_011+    1196113.9714827402
Rh001_043_011-    i_043    tia_h_in_001_011-    152446.63289477408
Rh001_044_011+    i_044    tia_h_in_001_011+    1189792.6169343942
Rh001_044_011-    i_044    tia_h_in_001_011-    259686.15732557568
Rh001_045_011+    i_045    tia_h_in_001_011+    1210646.6671559615
Rh001_045_011-    i_045    tia_h_in_001_011-    85982.27757007927
Rh001_046_011+    i_046    tia_h_in_001_011+    1199162.2346027293
Rh001_046_011-    i_046    tia_h_in_001_011-    238774.2200381138
Rh001_047_011+    i_047    tia_h_in_001_011+    67797.94774660612
Rh001_047_011-    i_047    tia_h_in_001_011-    1207091.4132740737
Rh001_048_011+    i_048    tia_h_in_001_011+    188522.20929642714
Rh001_048_011-    i_048    tia_h_in_001_011-    1189442.9562611424
Rh001_049_011+    i_049    tia_h_in_001_011+    1220822.5531786333
Rh001_049_011-    i_049    tia_h_in_001_011-    1014796.7638556177
Rh001_050_011+    i_050    tia_h_in_001_011+    84012.31358667882
Rh001_050_011-    i_050    tia_h_in_001_011-    1199889.1670533326
Rh001_051_011+    i_051    tia_h_in_001_011+    81028.20727462028
Rh001_051_011-    i_051    tia_h_in_001_011-    1207148.9967098157
Rh001_052_011+    i_052    tia_h_in_001_011+    81615.3019878155
Rh001_052_011-    i_052    tia_h_in_001_011-    1203376.2855601998
Rh001_053_011+    i_053    tia_h_in_001_011+    64192.04460659034
Rh001_053_011-    i_053    tia_h_in_001_011-    1190215.9114813237
Rh001_054_011+    i_054    tia_h_in_001_011+    266345.0126970063
Rh001_054_011-    i_054    tia_h_in_001_011-    1218686.2602184245
Rh001_055_011+    i_055    tia_h_in_001_011+    1181252.0947662692
Rh001_055_011-    i_055    tia_h_in_001_011-    83664.74281107892
Rh001_056_011+    i_056    tia_h_in_001_011+    72952.19985494259
Rh001_056_011-    i_056    tia_h_in_001_011-    1202062.1843857516
Rh001_057_011+    i_057    tia_h_in_001_011+    90216.16068791178
Rh001_057_011-    i_057    tia_h_in_001_011-    1218339.0812724505
Rh001_058_011+    i_058    tia_h_in_001_011+    228258.81216534358
Rh001_058_011-    i_058    tia_h_in_001_011-    1197239.4903176092
Rh001_059_011+    i_059    tia_h_in_001_011+    53813.81682523734
Rh001_059_011-    i_059    tia_h_in_001_011-    1197440.819856816
Rh001_060_011+    i_060    tia_h_in_001_011+    134450.7292547053
Rh001_060_011-    i_060    tia_h_in_001_011-    1201559.780172134
Rh001_061_011+    i_061    tia_h_in_001_011+    83940.58742824514
Rh001_061_011-    i_061    tia_h_in_001_011-    1199116.9184197832
Rh001_062_011+    i_062    tia_h_in_001_011+    217283.70724267457
Rh001_062_011-    i_062    tia_h_in_001_011-    1206787.829650878
Rh001_063_011+    i_063    tia_h_in_001_011+    45407.15573085015
Rh001_063_011-    i_063    tia_h_in_001_011-    1184478.4358348793
Rh001_064_011+    i_064    tia_h_in_001_011+    186341.8605851707
Rh001_064_011-    i_064    tia_h_in_001_011-    1214650.5308567253

* Neuron 12
Rh001_001_012+    i_001    tia_h_in_001_012+    1226036.871849852
Rh001_001_012-    i_001    tia_h_in_001_012-    61749.203495259266
Rh001_002_012+    i_002    tia_h_in_001_012+    254421.33857183185
Rh001_002_012-    i_002    tia_h_in_001_012-    1209263.6470815446
Rh001_003_012+    i_003    tia_h_in_001_012+    1193336.7287452824
Rh001_003_012-    i_003    tia_h_in_001_012-    63634.928895342215
Rh001_004_012+    i_004    tia_h_in_001_012+    49620.201557964276
Rh001_004_012-    i_004    tia_h_in_001_012-    1192962.261891149
Rh001_005_012+    i_005    tia_h_in_001_012+    68319.13942434969
Rh001_005_012-    i_005    tia_h_in_001_012-    1195206.5560608848
Rh001_006_012+    i_006    tia_h_in_001_012+    1203008.2280883982
Rh001_006_012-    i_006    tia_h_in_001_012-    266883.8351345649
Rh001_007_012+    i_007    tia_h_in_001_012+    134266.9785721228
Rh001_007_012-    i_007    tia_h_in_001_012-    1205969.5995339728
Rh001_008_012+    i_008    tia_h_in_001_012+    190149.90778246982
Rh001_008_012-    i_008    tia_h_in_001_012-    1187839.7791131365
Rh001_009_012+    i_009    tia_h_in_001_012+    107006.26102522161
Rh001_009_012-    i_009    tia_h_in_001_012-    1226988.4549469668
Rh001_010_012+    i_010    tia_h_in_001_012+    1191791.5880235399
Rh001_010_012-    i_010    tia_h_in_001_012-    73127.4176434589
Rh001_011_012+    i_011    tia_h_in_001_012+    1189886.3656101758
Rh001_011_012-    i_011    tia_h_in_001_012-    555965.1812104167
Rh001_012_012+    i_012    tia_h_in_001_012+    1201193.0530663193
Rh001_012_012-    i_012    tia_h_in_001_012-    94570.05039064311
Rh001_013_012+    i_013    tia_h_in_001_012+    95274.85110828659
Rh001_013_012-    i_013    tia_h_in_001_012-    1194155.4974679847
Rh001_014_012+    i_014    tia_h_in_001_012+    47943.11434514576
Rh001_014_012-    i_014    tia_h_in_001_012-    1204207.9456014212
Rh001_015_012+    i_015    tia_h_in_001_012+    78620.23541793112
Rh001_015_012-    i_015    tia_h_in_001_012-    1199384.639752062
Rh001_016_012+    i_016    tia_h_in_001_012+    104213.18254044277
Rh001_016_012-    i_016    tia_h_in_001_012-    1185648.9075514576
Rh001_017_012+    i_017    tia_h_in_001_012+    1204257.7962760378
Rh001_017_012-    i_017    tia_h_in_001_012-    272500.0999351388
Rh001_018_012+    i_018    tia_h_in_001_012+    46061.987527189915
Rh001_018_012-    i_018    tia_h_in_001_012-    1202727.1847995135
Rh001_019_012+    i_019    tia_h_in_001_012+    92280.26130360799
Rh001_019_012-    i_019    tia_h_in_001_012-    1202954.9507423271
Rh001_020_012+    i_020    tia_h_in_001_012+    1211991.4466451304
Rh001_020_012-    i_020    tia_h_in_001_012-    48972.056659330694
Rh001_021_012+    i_021    tia_h_in_001_012+    218257.53689900308
Rh001_021_012-    i_021    tia_h_in_001_012-    1203687.9017574547
Rh001_022_012+    i_022    tia_h_in_001_012+    1202006.3818609393
Rh001_022_012-    i_022    tia_h_in_001_012-    288586.1537752873
Rh001_023_012+    i_023    tia_h_in_001_012+    47118.88338632002
Rh001_023_012-    i_023    tia_h_in_001_012-    1178106.78886009
Rh001_024_012+    i_024    tia_h_in_001_012+    280829.1470309589
Rh001_024_012-    i_024    tia_h_in_001_012-    1208076.7996916901
Rh001_025_012+    i_025    tia_h_in_001_012+    1193739.5817020836
Rh001_025_012-    i_025    tia_h_in_001_012-    96182.00431149003
Rh001_026_012+    i_026    tia_h_in_001_012+    96237.75173095806
Rh001_026_012-    i_026    tia_h_in_001_012-    1188065.1337075466
Rh001_027_012+    i_027    tia_h_in_001_012+    43512.30577629223
Rh001_027_012-    i_027    tia_h_in_001_012-    1214024.632155025
Rh001_028_012+    i_028    tia_h_in_001_012+    65331.37446291168
Rh001_028_012-    i_028    tia_h_in_001_012-    1204567.195981981
Rh001_029_012+    i_029    tia_h_in_001_012+    234380.67208052005
Rh001_029_012-    i_029    tia_h_in_001_012-    1184151.9540949736
Rh001_030_012+    i_030    tia_h_in_001_012+    286943.24958040525
Rh001_030_012-    i_030    tia_h_in_001_012-    1196453.535997841
Rh001_031_012+    i_031    tia_h_in_001_012+    49542.25792812123
Rh001_031_012-    i_031    tia_h_in_001_012-    1202187.9943046188
Rh001_032_012+    i_032    tia_h_in_001_012+    30464.82337480282
Rh001_032_012-    i_032    tia_h_in_001_012-    1206960.345605833
Rh001_033_012+    i_033    tia_h_in_001_012+    50495.27195691368
Rh001_033_012-    i_033    tia_h_in_001_012-    1206890.7762204173
Rh001_034_012+    i_034    tia_h_in_001_012+    148810.744899411
Rh001_034_012-    i_034    tia_h_in_001_012-    1203103.7018474478
Rh001_035_012+    i_035    tia_h_in_001_012+    67239.28456266536
Rh001_035_012-    i_035    tia_h_in_001_012-    1198437.3219839244
Rh001_036_012+    i_036    tia_h_in_001_012+    118613.29174878585
Rh001_036_012-    i_036    tia_h_in_001_012-    1211217.206512051
Rh001_037_012+    i_037    tia_h_in_001_012+    100720.77526661761
Rh001_037_012-    i_037    tia_h_in_001_012-    1193853.8626032493
Rh001_038_012+    i_038    tia_h_in_001_012+    107213.14685795641
Rh001_038_012-    i_038    tia_h_in_001_012-    1202384.0131752202
Rh001_039_012+    i_039    tia_h_in_001_012+    72905.64849426915
Rh001_039_012-    i_039    tia_h_in_001_012-    1190359.3135039129
Rh001_040_012+    i_040    tia_h_in_001_012+    1201678.7717730328
Rh001_040_012-    i_040    tia_h_in_001_012-    238066.78185518167
Rh001_041_012+    i_041    tia_h_in_001_012+    40617.8000272474
Rh001_041_012-    i_041    tia_h_in_001_012-    1196020.69764616
Rh001_042_012+    i_042    tia_h_in_001_012+    66370.1690167202
Rh001_042_012-    i_042    tia_h_in_001_012-    1186366.9888671471
Rh001_043_012+    i_043    tia_h_in_001_012+    129679.6307171327
Rh001_043_012-    i_043    tia_h_in_001_012-    1198419.5821853427
Rh001_044_012+    i_044    tia_h_in_001_012+    69218.14310597682
Rh001_044_012-    i_044    tia_h_in_001_012-    1192725.6231753868
Rh001_045_012+    i_045    tia_h_in_001_012+    1211174.4925921874
Rh001_045_012-    i_045    tia_h_in_001_012-    189938.2669348269
Rh001_046_012+    i_046    tia_h_in_001_012+    1203448.4729590984
Rh001_046_012-    i_046    tia_h_in_001_012-    133570.8522935707
Rh001_047_012+    i_047    tia_h_in_001_012+    86160.4967645649
Rh001_047_012-    i_047    tia_h_in_001_012-    1206915.9453261753
Rh001_048_012+    i_048    tia_h_in_001_012+    1185516.8995090646
Rh001_048_012-    i_048    tia_h_in_001_012-    121825.60505707705
Rh001_049_012+    i_049    tia_h_in_001_012+    49461.001229949616
Rh001_049_012-    i_049    tia_h_in_001_012-    1209877.8243041951
Rh001_050_012+    i_050    tia_h_in_001_012+    52844.33238474716
Rh001_050_012-    i_050    tia_h_in_001_012-    1201689.3856889354
Rh001_051_012+    i_051    tia_h_in_001_012+    273642.3480443491
Rh001_051_012-    i_051    tia_h_in_001_012-    1203967.067517368
Rh001_052_012+    i_052    tia_h_in_001_012+    90520.59300761923
Rh001_052_012-    i_052    tia_h_in_001_012-    1200009.5270171685
Rh001_053_012+    i_053    tia_h_in_001_012+    35256.95518498427
Rh001_053_012-    i_053    tia_h_in_001_012-    1189076.7616554825
Rh001_054_012+    i_054    tia_h_in_001_012+    76729.28794456532
Rh001_054_012-    i_054    tia_h_in_001_012-    1215086.937323075
Rh001_055_012+    i_055    tia_h_in_001_012+    1199044.675385433
Rh001_055_012-    i_055    tia_h_in_001_012-    165938.88310053977
Rh001_056_012+    i_056    tia_h_in_001_012+    131701.84363099543
Rh001_056_012-    i_056    tia_h_in_001_012-    1196482.9115766468
Rh001_057_012+    i_057    tia_h_in_001_012+    1205882.9473644132
Rh001_057_012-    i_057    tia_h_in_001_012-    151118.11132011475
Rh001_058_012+    i_058    tia_h_in_001_012+    101600.08132562488
Rh001_058_012-    i_058    tia_h_in_001_012-    1209273.1997725223
Rh001_059_012+    i_059    tia_h_in_001_012+    1205768.2948424416
Rh001_059_012-    i_059    tia_h_in_001_012-    221478.2371403517
Rh001_060_012+    i_060    tia_h_in_001_012+    1197275.0024698083
Rh001_060_012-    i_060    tia_h_in_001_012-    177293.947941562
Rh001_061_012+    i_061    tia_h_in_001_012+    76807.82886916852
Rh001_061_012-    i_061    tia_h_in_001_012-    1205530.974823422
Rh001_062_012+    i_062    tia_h_in_001_012+    1201552.1752138948
Rh001_062_012-    i_062    tia_h_in_001_012-    132634.868249281
Rh001_063_012+    i_063    tia_h_in_001_012+    1205342.6574237496
Rh001_063_012-    i_063    tia_h_in_001_012-    89386.84031280316
Rh001_064_012+    i_064    tia_h_in_001_012+    1215929.4289668973
Rh001_064_012-    i_064    tia_h_in_001_012-    581927.8491738752

* Neuron 13
Rh001_001_013+    i_001    tia_h_in_001_013+    1177308.9633597091
Rh001_001_013-    i_001    tia_h_in_001_013-    26916.756912159788
Rh001_002_013+    i_002    tia_h_in_001_013+    1195355.50735884
Rh001_002_013-    i_002    tia_h_in_001_013-    25830.421910070156
Rh001_003_013+    i_003    tia_h_in_001_013+    1190279.3017768415
Rh001_003_013-    i_003    tia_h_in_001_013-    78858.76820818974
Rh001_004_013+    i_004    tia_h_in_001_013+    1212227.695098559
Rh001_004_013-    i_004    tia_h_in_001_013-    95662.94311765974
Rh001_005_013+    i_005    tia_h_in_001_013+    1200682.3670506305
Rh001_005_013-    i_005    tia_h_in_001_013-    253258.56833696133
Rh001_006_013+    i_006    tia_h_in_001_013+    61371.869312215764
Rh001_006_013-    i_006    tia_h_in_001_013-    1203984.2974286904
Rh001_007_013+    i_007    tia_h_in_001_013+    1209594.2400265737
Rh001_007_013-    i_007    tia_h_in_001_013-    1011606.3664025472
Rh001_008_013+    i_008    tia_h_in_001_013+    66653.92929940486
Rh001_008_013-    i_008    tia_h_in_001_013-    1198573.3765211515
Rh001_009_013+    i_009    tia_h_in_001_013+    81932.61586228604
Rh001_009_013-    i_009    tia_h_in_001_013-    1196462.5878859686
Rh001_010_013+    i_010    tia_h_in_001_013+    93022.19732248783
Rh001_010_013-    i_010    tia_h_in_001_013-    1197695.060819173
Rh001_011_013+    i_011    tia_h_in_001_013+    49552.10822585455
Rh001_011_013-    i_011    tia_h_in_001_013-    1212662.8211893719
Rh001_012_013+    i_012    tia_h_in_001_013+    1195172.859691459
Rh001_012_013-    i_012    tia_h_in_001_013-    504517.02313150984
Rh001_013_013+    i_013    tia_h_in_001_013+    168569.70908311068
Rh001_013_013-    i_013    tia_h_in_001_013-    1193441.044615784
Rh001_014_013+    i_014    tia_h_in_001_013+    1191881.4212905637
Rh001_014_013-    i_014    tia_h_in_001_013-    434620.67823607335
Rh001_015_013+    i_015    tia_h_in_001_013+    104882.53053661472
Rh001_015_013-    i_015    tia_h_in_001_013-    1207350.1967267164
Rh001_016_013+    i_016    tia_h_in_001_013+    90363.9539409886
Rh001_016_013-    i_016    tia_h_in_001_013-    1194625.4173828051
Rh001_017_013+    i_017    tia_h_in_001_013+    25346.322386927575
Rh001_017_013-    i_017    tia_h_in_001_013-    1206883.2870958743
Rh001_018_013+    i_018    tia_h_in_001_013+    42537.74410243981
Rh001_018_013-    i_018    tia_h_in_001_013-    1202957.4351733583
Rh001_019_013+    i_019    tia_h_in_001_013+    47283.057718530006
Rh001_019_013-    i_019    tia_h_in_001_013-    1199733.835001172
Rh001_020_013+    i_020    tia_h_in_001_013+    110920.76946112675
Rh001_020_013-    i_020    tia_h_in_001_013-    1191275.443910109
Rh001_021_013+    i_021    tia_h_in_001_013+    575470.1924927405
Rh001_021_013-    i_021    tia_h_in_001_013-    1196278.2126819054
Rh001_022_013+    i_022    tia_h_in_001_013+    1210634.8419519835
Rh001_022_013-    i_022    tia_h_in_001_013-    598071.8007444448
Rh001_023_013+    i_023    tia_h_in_001_013+    1202830.4787752565
Rh001_023_013-    i_023    tia_h_in_001_013-    165314.03996282865
Rh001_024_013+    i_024    tia_h_in_001_013+    1199547.9592986212
Rh001_024_013-    i_024    tia_h_in_001_013-    59432.52259216932
Rh001_025_013+    i_025    tia_h_in_001_013+    52113.12352318112
Rh001_025_013-    i_025    tia_h_in_001_013-    1194801.930105261
Rh001_026_013+    i_026    tia_h_in_001_013+    73300.72010572653
Rh001_026_013-    i_026    tia_h_in_001_013-    1199403.6476908142
Rh001_027_013+    i_027    tia_h_in_001_013+    59736.840948585545
Rh001_027_013-    i_027    tia_h_in_001_013-    1192284.8324750033
Rh001_028_013+    i_028    tia_h_in_001_013+    68673.23246145509
Rh001_028_013-    i_028    tia_h_in_001_013-    1196262.7816477553
Rh001_029_013+    i_029    tia_h_in_001_013+    1204340.674161749
Rh001_029_013-    i_029    tia_h_in_001_013-    79674.4607145986
Rh001_030_013+    i_030    tia_h_in_001_013+    73161.30153857052
Rh001_030_013-    i_030    tia_h_in_001_013-    1198574.4357729778
Rh001_031_013+    i_031    tia_h_in_001_013+    328898.83071001974
Rh001_031_013-    i_031    tia_h_in_001_013-    1205311.1898812482
Rh001_032_013+    i_032    tia_h_in_001_013+    78609.3210772291
Rh001_032_013-    i_032    tia_h_in_001_013-    1225592.7679517136
Rh001_033_013+    i_033    tia_h_in_001_013+    410891.1258313932
Rh001_033_013-    i_033    tia_h_in_001_013-    1196435.1719524025
Rh001_034_013+    i_034    tia_h_in_001_013+    1202749.1414945535
Rh001_034_013-    i_034    tia_h_in_001_013-    1160096.9659110797
Rh001_035_013+    i_035    tia_h_in_001_013+    173482.8399427413
Rh001_035_013-    i_035    tia_h_in_001_013-    1208602.7696324375
Rh001_036_013+    i_036    tia_h_in_001_013+    133093.3765364676
Rh001_036_013-    i_036    tia_h_in_001_013-    1199790.9719242232
Rh001_037_013+    i_037    tia_h_in_001_013+    38697.06971478538
Rh001_037_013-    i_037    tia_h_in_001_013-    1199102.2398334132
Rh001_038_013+    i_038    tia_h_in_001_013+    536658.7446959482
Rh001_038_013-    i_038    tia_h_in_001_013-    1190618.015755214
Rh001_039_013+    i_039    tia_h_in_001_013+    118739.00213941497
Rh001_039_013-    i_039    tia_h_in_001_013-    1212522.4053297827
Rh001_040_013+    i_040    tia_h_in_001_013+    1216034.989041206
Rh001_040_013-    i_040    tia_h_in_001_013-    628457.1830142026
Rh001_041_013+    i_041    tia_h_in_001_013+    1195023.1831451969
Rh001_041_013-    i_041    tia_h_in_001_013-    1206533.8746936624
Rh001_042_013+    i_042    tia_h_in_001_013+    90555.33297578107
Rh001_042_013-    i_042    tia_h_in_001_013-    1179822.9571741968
Rh001_043_013+    i_043    tia_h_in_001_013+    130416.96151492096
Rh001_043_013-    i_043    tia_h_in_001_013-    1197020.9000490222
Rh001_044_013+    i_044    tia_h_in_001_013+    114872.02512030149
Rh001_044_013-    i_044    tia_h_in_001_013-    1212885.3930966817
Rh001_045_013+    i_045    tia_h_in_001_013+    34498.73926015158
Rh001_045_013-    i_045    tia_h_in_001_013-    1206380.8560297256
Rh001_046_013+    i_046    tia_h_in_001_013+    39037.65971106016
Rh001_046_013-    i_046    tia_h_in_001_013-    1186591.8665808304
Rh001_047_013+    i_047    tia_h_in_001_013+    50971.27549352147
Rh001_047_013-    i_047    tia_h_in_001_013-    1203096.278444395
Rh001_048_013+    i_048    tia_h_in_001_013+    238954.59753414293
Rh001_048_013-    i_048    tia_h_in_001_013-    1198436.7431316036
Rh001_049_013+    i_049    tia_h_in_001_013+    828364.5905158968
Rh001_049_013-    i_049    tia_h_in_001_013-    1215680.8270069456
Rh001_050_013+    i_050    tia_h_in_001_013+    176179.2615085833
Rh001_050_013-    i_050    tia_h_in_001_013-    1185079.2141577075
Rh001_051_013+    i_051    tia_h_in_001_013+    111621.86602783404
Rh001_051_013-    i_051    tia_h_in_001_013-    1204401.6415181877
Rh001_052_013+    i_052    tia_h_in_001_013+    1201725.8359959049
Rh001_052_013-    i_052    tia_h_in_001_013-    470503.28608951136
Rh001_053_013+    i_053    tia_h_in_001_013+    1211983.6222134756
Rh001_053_013-    i_053    tia_h_in_001_013-    699509.8546240554
Rh001_054_013+    i_054    tia_h_in_001_013+    64713.26025522371
Rh001_054_013-    i_054    tia_h_in_001_013-    1187304.6626838585
Rh001_055_013+    i_055    tia_h_in_001_013+    81200.9097668717
Rh001_055_013-    i_055    tia_h_in_001_013-    1185709.0948532207
Rh001_056_013+    i_056    tia_h_in_001_013+    105346.66414980637
Rh001_056_013-    i_056    tia_h_in_001_013-    1190727.072600911
Rh001_057_013+    i_057    tia_h_in_001_013+    55533.5784477653
Rh001_057_013-    i_057    tia_h_in_001_013-    1204210.3860930272
Rh001_058_013+    i_058    tia_h_in_001_013+    301017.69347983133
Rh001_058_013-    i_058    tia_h_in_001_013-    1190120.3233325132
Rh001_059_013+    i_059    tia_h_in_001_013+    260497.97466534836
Rh001_059_013-    i_059    tia_h_in_001_013-    1193723.9104708587
Rh001_060_013+    i_060    tia_h_in_001_013+    70831.85886801693
Rh001_060_013-    i_060    tia_h_in_001_013-    1189834.0380586006
Rh001_061_013+    i_061    tia_h_in_001_013+    167693.11269889676
Rh001_061_013-    i_061    tia_h_in_001_013-    1197273.9922823883
Rh001_062_013+    i_062    tia_h_in_001_013+    317539.97896751185
Rh001_062_013-    i_062    tia_h_in_001_013-    1184365.2247871503
Rh001_063_013+    i_063    tia_h_in_001_013+    1200688.3157454592
Rh001_063_013-    i_063    tia_h_in_001_013-    175795.0130319518
Rh001_064_013+    i_064    tia_h_in_001_013+    59646.09098081393
Rh001_064_013-    i_064    tia_h_in_001_013-    1187685.3494343816

* Neuron 14
Rh001_001_014+    i_001    tia_h_in_001_014+    1202317.7158355345
Rh001_001_014-    i_001    tia_h_in_001_014-    423469.5414650479
Rh001_002_014+    i_002    tia_h_in_001_014+    197041.3670016536
Rh001_002_014-    i_002    tia_h_in_001_014-    1195438.5198015058
Rh001_003_014+    i_003    tia_h_in_001_014+    131720.3086458252
Rh001_003_014-    i_003    tia_h_in_001_014-    1170176.5583881137
Rh001_004_014+    i_004    tia_h_in_001_014+    850877.2843111363
Rh001_004_014-    i_004    tia_h_in_001_014-    1209996.8188877858
Rh001_005_014+    i_005    tia_h_in_001_014+    112854.1898219527
Rh001_005_014-    i_005    tia_h_in_001_014-    1202938.9693630177
Rh001_006_014+    i_006    tia_h_in_001_014+    1206192.0579338134
Rh001_006_014-    i_006    tia_h_in_001_014-    208914.69213328205
Rh001_007_014+    i_007    tia_h_in_001_014+    1192572.9177781288
Rh001_007_014-    i_007    tia_h_in_001_014-    424249.21586242085
Rh001_008_014+    i_008    tia_h_in_001_014+    1201520.3072648689
Rh001_008_014-    i_008    tia_h_in_001_014-    220372.39170567636
Rh001_009_014+    i_009    tia_h_in_001_014+    360726.7316411323
Rh001_009_014-    i_009    tia_h_in_001_014-    1202237.1285876145
Rh001_010_014+    i_010    tia_h_in_001_014+    475427.00218272867
Rh001_010_014-    i_010    tia_h_in_001_014-    1204002.5050484992
Rh001_011_014+    i_011    tia_h_in_001_014+    139433.14863988588
Rh001_011_014-    i_011    tia_h_in_001_014-    1205136.9301559944
Rh001_012_014+    i_012    tia_h_in_001_014+    255033.12439588326
Rh001_012_014-    i_012    tia_h_in_001_014-    1198102.1933129006
Rh001_013_014+    i_013    tia_h_in_001_014+    99393.05848709698
Rh001_013_014-    i_013    tia_h_in_001_014-    1203622.4169289852
Rh001_014_014+    i_014    tia_h_in_001_014+    71227.34566100402
Rh001_014_014-    i_014    tia_h_in_001_014-    1191590.7647833768
Rh001_015_014+    i_015    tia_h_in_001_014+    112714.76440418158
Rh001_015_014-    i_015    tia_h_in_001_014-    1190198.73715083
Rh001_016_014+    i_016    tia_h_in_001_014+    770295.8132252914
Rh001_016_014-    i_016    tia_h_in_001_014-    1214684.9925458143
Rh001_017_014+    i_017    tia_h_in_001_014+    1206050.8240911986
Rh001_017_014-    i_017    tia_h_in_001_014-    269611.8896288248
Rh001_018_014+    i_018    tia_h_in_001_014+    106684.51866540892
Rh001_018_014-    i_018    tia_h_in_001_014-    1189802.3252931517
Rh001_019_014+    i_019    tia_h_in_001_014+    550833.7007219703
Rh001_019_014-    i_019    tia_h_in_001_014-    1215688.7811543904
Rh001_020_014+    i_020    tia_h_in_001_014+    95919.33879771281
Rh001_020_014-    i_020    tia_h_in_001_014-    1197304.2088727658
Rh001_021_014+    i_021    tia_h_in_001_014+    88470.15014076636
Rh001_021_014-    i_021    tia_h_in_001_014-    1182769.2438925162
Rh001_022_014+    i_022    tia_h_in_001_014+    110291.56327912441
Rh001_022_014-    i_022    tia_h_in_001_014-    1209017.227572735
Rh001_023_014+    i_023    tia_h_in_001_014+    71578.51339421733
Rh001_023_014-    i_023    tia_h_in_001_014-    1198437.965403959
Rh001_024_014+    i_024    tia_h_in_001_014+    74062.04144400214
Rh001_024_014-    i_024    tia_h_in_001_014-    1182489.7036040304
Rh001_025_014+    i_025    tia_h_in_001_014+    126749.0386739939
Rh001_025_014-    i_025    tia_h_in_001_014-    1198397.4847741723
Rh001_026_014+    i_026    tia_h_in_001_014+    1212435.7631726426
Rh001_026_014-    i_026    tia_h_in_001_014-    590628.6500594879
Rh001_027_014+    i_027    tia_h_in_001_014+    69992.39981718925
Rh001_027_014-    i_027    tia_h_in_001_014-    1199872.7705507723
Rh001_028_014+    i_028    tia_h_in_001_014+    540725.7473834886
Rh001_028_014-    i_028    tia_h_in_001_014-    1184985.0295842695
Rh001_029_014+    i_029    tia_h_in_001_014+    1124975.6976316157
Rh001_029_014-    i_029    tia_h_in_001_014-    1195501.6444599098
Rh001_030_014+    i_030    tia_h_in_001_014+    75398.8573466484
Rh001_030_014-    i_030    tia_h_in_001_014-    1194018.9554577908
Rh001_031_014+    i_031    tia_h_in_001_014+    80442.73134947305
Rh001_031_014-    i_031    tia_h_in_001_014-    1186434.8410439496
Rh001_032_014+    i_032    tia_h_in_001_014+    125609.11665368766
Rh001_032_014-    i_032    tia_h_in_001_014-    1213279.5498537845
Rh001_033_014+    i_033    tia_h_in_001_014+    174548.19882241398
Rh001_033_014-    i_033    tia_h_in_001_014-    1218125.5955664688
Rh001_034_014+    i_034    tia_h_in_001_014+    1202360.5445260007
Rh001_034_014-    i_034    tia_h_in_001_014-    333276.4384113674
Rh001_035_014+    i_035    tia_h_in_001_014+    204242.11562636044
Rh001_035_014-    i_035    tia_h_in_001_014-    1198767.5280454087
Rh001_036_014+    i_036    tia_h_in_001_014+    66943.28398512429
Rh001_036_014-    i_036    tia_h_in_001_014-    1211348.3506289923
Rh001_037_014+    i_037    tia_h_in_001_014+    128672.04028297712
Rh001_037_014-    i_037    tia_h_in_001_014-    1197062.3944210792
Rh001_038_014+    i_038    tia_h_in_001_014+    158144.53243487707
Rh001_038_014-    i_038    tia_h_in_001_014-    1215135.0780221866
Rh001_039_014+    i_039    tia_h_in_001_014+    297249.56689439365
Rh001_039_014-    i_039    tia_h_in_001_014-    1202447.489252084
Rh001_040_014+    i_040    tia_h_in_001_014+    344116.85881619394
Rh001_040_014-    i_040    tia_h_in_001_014-    1211566.7487913545
Rh001_041_014+    i_041    tia_h_in_001_014+    93517.2357286041
Rh001_041_014-    i_041    tia_h_in_001_014-    1198255.4294182074
Rh001_042_014+    i_042    tia_h_in_001_014+    167841.052210831
Rh001_042_014-    i_042    tia_h_in_001_014-    1199926.425206783
Rh001_043_014+    i_043    tia_h_in_001_014+    88925.68795100528
Rh001_043_014-    i_043    tia_h_in_001_014-    1195093.0901679925
Rh001_044_014+    i_044    tia_h_in_001_014+    229972.94478992085
Rh001_044_014-    i_044    tia_h_in_001_014-    1194471.666760108
Rh001_045_014+    i_045    tia_h_in_001_014+    100086.42441084699
Rh001_045_014-    i_045    tia_h_in_001_014-    1181876.260746998
Rh001_046_014+    i_046    tia_h_in_001_014+    106508.97546463834
Rh001_046_014-    i_046    tia_h_in_001_014-    1201427.9279833534
Rh001_047_014+    i_047    tia_h_in_001_014+    144029.62825340877
Rh001_047_014-    i_047    tia_h_in_001_014-    1200401.7208544377
Rh001_048_014+    i_048    tia_h_in_001_014+    80717.68828401073
Rh001_048_014-    i_048    tia_h_in_001_014-    1196324.5695144888
Rh001_049_014+    i_049    tia_h_in_001_014+    93872.28988005061
Rh001_049_014-    i_049    tia_h_in_001_014-    1208564.423953856
Rh001_050_014+    i_050    tia_h_in_001_014+    74147.26830207279
Rh001_050_014-    i_050    tia_h_in_001_014-    1202013.3788502424
Rh001_051_014+    i_051    tia_h_in_001_014+    84183.00568930939
Rh001_051_014-    i_051    tia_h_in_001_014-    1207483.4300832043
Rh001_052_014+    i_052    tia_h_in_001_014+    337168.3517049982
Rh001_052_014-    i_052    tia_h_in_001_014-    1202206.4969903515
Rh001_053_014+    i_053    tia_h_in_001_014+    1205285.8325799992
Rh001_053_014-    i_053    tia_h_in_001_014-    274421.5059273569
Rh001_054_014+    i_054    tia_h_in_001_014+    146112.87406963424
Rh001_054_014-    i_054    tia_h_in_001_014-    1197840.733770366
Rh001_055_014+    i_055    tia_h_in_001_014+    175434.34076371993
Rh001_055_014-    i_055    tia_h_in_001_014-    1203278.9548637941
Rh001_056_014+    i_056    tia_h_in_001_014+    249266.65835577392
Rh001_056_014-    i_056    tia_h_in_001_014-    1197946.2210930435
Rh001_057_014+    i_057    tia_h_in_001_014+    300021.3292596241
Rh001_057_014-    i_057    tia_h_in_001_014-    1226429.120646019
Rh001_058_014+    i_058    tia_h_in_001_014+    188046.36092904818
Rh001_058_014-    i_058    tia_h_in_001_014-    1205392.6041247854
Rh001_059_014+    i_059    tia_h_in_001_014+    86771.58949491334
Rh001_059_014-    i_059    tia_h_in_001_014-    1193263.9928297945
Rh001_060_014+    i_060    tia_h_in_001_014+    124186.67272459225
Rh001_060_014-    i_060    tia_h_in_001_014-    1189754.6393137556
Rh001_061_014+    i_061    tia_h_in_001_014+    375294.71005721635
Rh001_061_014-    i_061    tia_h_in_001_014-    1194341.8090324446
Rh001_062_014+    i_062    tia_h_in_001_014+    559913.6617344237
Rh001_062_014-    i_062    tia_h_in_001_014-    1180437.2511055693
Rh001_063_014+    i_063    tia_h_in_001_014+    251526.56630069765
Rh001_063_014-    i_063    tia_h_in_001_014-    1190894.8265461926
Rh001_064_014+    i_064    tia_h_in_001_014+    424806.92085503327
Rh001_064_014-    i_064    tia_h_in_001_014-    1207103.0953638353

* Neuron 15
Rh001_001_015+    i_001    tia_h_in_001_015+    67860.28737035462
Rh001_001_015-    i_001    tia_h_in_001_015-    1206511.5681555553
Rh001_002_015+    i_002    tia_h_in_001_015+    88665.74262149211
Rh001_002_015-    i_002    tia_h_in_001_015-    1207490.634219297
Rh001_003_015+    i_003    tia_h_in_001_015+    67399.46577323765
Rh001_003_015-    i_003    tia_h_in_001_015-    1211239.920079641
Rh001_004_015+    i_004    tia_h_in_001_015+    149755.0615071737
Rh001_004_015-    i_004    tia_h_in_001_015-    1195784.0757427288
Rh001_005_015+    i_005    tia_h_in_001_015+    121378.67771949843
Rh001_005_015-    i_005    tia_h_in_001_015-    1192478.81391973
Rh001_006_015+    i_006    tia_h_in_001_015+    103439.95605779054
Rh001_006_015-    i_006    tia_h_in_001_015-    1199846.7061248245
Rh001_007_015+    i_007    tia_h_in_001_015+    1189435.6366970937
Rh001_007_015-    i_007    tia_h_in_001_015-    281102.66304013535
Rh001_008_015+    i_008    tia_h_in_001_015+    134909.4995976199
Rh001_008_015-    i_008    tia_h_in_001_015-    1195640.0152984937
Rh001_009_015+    i_009    tia_h_in_001_015+    162228.81371360586
Rh001_009_015-    i_009    tia_h_in_001_015-    1200076.0043586337
Rh001_010_015+    i_010    tia_h_in_001_015+    702263.557920113
Rh001_010_015-    i_010    tia_h_in_001_015-    1201318.9568919889
Rh001_011_015+    i_011    tia_h_in_001_015+    1194380.602875384
Rh001_011_015-    i_011    tia_h_in_001_015-    488250.30733795604
Rh001_012_015+    i_012    tia_h_in_001_015+    68405.37528781094
Rh001_012_015-    i_012    tia_h_in_001_015-    1197191.8983192828
Rh001_013_015+    i_013    tia_h_in_001_015+    72519.88693576798
Rh001_013_015-    i_013    tia_h_in_001_015-    1208259.6304139735
Rh001_014_015+    i_014    tia_h_in_001_015+    93418.89498209287
Rh001_014_015-    i_014    tia_h_in_001_015-    1199097.8659451483
Rh001_015_015+    i_015    tia_h_in_001_015+    66706.69126202777
Rh001_015_015-    i_015    tia_h_in_001_015-    1200179.0919265626
Rh001_016_015+    i_016    tia_h_in_001_015+    325465.52369199
Rh001_016_015-    i_016    tia_h_in_001_015-    1189723.9299217372
Rh001_017_015+    i_017    tia_h_in_001_015+    195379.5102563779
Rh001_017_015-    i_017    tia_h_in_001_015-    1211195.2136422433
Rh001_018_015+    i_018    tia_h_in_001_015+    100315.53912608148
Rh001_018_015-    i_018    tia_h_in_001_015-    1214755.2366208786
Rh001_019_015+    i_019    tia_h_in_001_015+    193751.1035132903
Rh001_019_015-    i_019    tia_h_in_001_015-    1211597.3370201655
Rh001_020_015+    i_020    tia_h_in_001_015+    209319.13661583044
Rh001_020_015-    i_020    tia_h_in_001_015-    1200887.3873588364
Rh001_021_015+    i_021    tia_h_in_001_015+    1192054.5984592503
Rh001_021_015-    i_021    tia_h_in_001_015-    400397.71968533524
Rh001_022_015+    i_022    tia_h_in_001_015+    112887.78950759809
Rh001_022_015-    i_022    tia_h_in_001_015-    1205333.0219135548
Rh001_023_015+    i_023    tia_h_in_001_015+    857433.8691069495
Rh001_023_015-    i_023    tia_h_in_001_015-    1196326.21813926
Rh001_024_015+    i_024    tia_h_in_001_015+    140335.6559111799
Rh001_024_015-    i_024    tia_h_in_001_015-    1209298.6997484975
Rh001_025_015+    i_025    tia_h_in_001_015+    65336.26962457402
Rh001_025_015-    i_025    tia_h_in_001_015-    1194120.9464027476
Rh001_026_015+    i_026    tia_h_in_001_015+    259068.80531572897
Rh001_026_015-    i_026    tia_h_in_001_015-    1202528.129025811
Rh001_027_015+    i_027    tia_h_in_001_015+    262484.11831021786
Rh001_027_015-    i_027    tia_h_in_001_015-    1184861.729036264
Rh001_028_015+    i_028    tia_h_in_001_015+    83005.8507808319
Rh001_028_015-    i_028    tia_h_in_001_015-    1206557.8136432078
Rh001_029_015+    i_029    tia_h_in_001_015+    299705.90221313393
Rh001_029_015-    i_029    tia_h_in_001_015-    1196593.338970442
Rh001_030_015+    i_030    tia_h_in_001_015+    181578.09121970867
Rh001_030_015-    i_030    tia_h_in_001_015-    1197094.627794753
Rh001_031_015+    i_031    tia_h_in_001_015+    65704.0690502901
Rh001_031_015-    i_031    tia_h_in_001_015-    1203796.898286233
Rh001_032_015+    i_032    tia_h_in_001_015+    337040.35144008824
Rh001_032_015-    i_032    tia_h_in_001_015-    1193126.1164731078
Rh001_033_015+    i_033    tia_h_in_001_015+    1200497.5092116985
Rh001_033_015-    i_033    tia_h_in_001_015-    679886.2669060911
Rh001_034_015+    i_034    tia_h_in_001_015+    641311.5249464528
Rh001_034_015-    i_034    tia_h_in_001_015-    1190547.5208927712
Rh001_035_015+    i_035    tia_h_in_001_015+    243017.10785122417
Rh001_035_015-    i_035    tia_h_in_001_015-    1204758.7704026774
Rh001_036_015+    i_036    tia_h_in_001_015+    423626.37626338727
Rh001_036_015-    i_036    tia_h_in_001_015-    1184291.4823166074
Rh001_037_015+    i_037    tia_h_in_001_015+    507504.0374335114
Rh001_037_015-    i_037    tia_h_in_001_015-    1201881.8917114078
Rh001_038_015+    i_038    tia_h_in_001_015+    100540.60476807664
Rh001_038_015-    i_038    tia_h_in_001_015-    1200584.1176402501
Rh001_039_015+    i_039    tia_h_in_001_015+    125524.15836621156
Rh001_039_015-    i_039    tia_h_in_001_015-    1212208.0535763472
Rh001_040_015+    i_040    tia_h_in_001_015+    268600.4727225007
Rh001_040_015-    i_040    tia_h_in_001_015-    1194177.8305988135
Rh001_041_015+    i_041    tia_h_in_001_015+    1191001.4579689028
Rh001_041_015-    i_041    tia_h_in_001_015-    522143.3226908582
Rh001_042_015+    i_042    tia_h_in_001_015+    269390.754080323
Rh001_042_015-    i_042    tia_h_in_001_015-    1192041.3401237703
Rh001_043_015+    i_043    tia_h_in_001_015+    343738.71149982064
Rh001_043_015-    i_043    tia_h_in_001_015-    1197670.3450924144
Rh001_044_015+    i_044    tia_h_in_001_015+    273397.3046945038
Rh001_044_015-    i_044    tia_h_in_001_015-    1211053.0110281368
Rh001_045_015+    i_045    tia_h_in_001_015+    1210234.461144815
Rh001_045_015-    i_045    tia_h_in_001_015-    320064.18851280457
Rh001_046_015+    i_046    tia_h_in_001_015+    120018.60496815413
Rh001_046_015-    i_046    tia_h_in_001_015-    1199447.1806875463
Rh001_047_015+    i_047    tia_h_in_001_015+    1193094.5204147075
Rh001_047_015-    i_047    tia_h_in_001_015-    593141.2659714078
Rh001_048_015+    i_048    tia_h_in_001_015+    1194407.043755412
Rh001_048_015-    i_048    tia_h_in_001_015-    474972.10649888037
Rh001_049_015+    i_049    tia_h_in_001_015+    1200646.7849172107
Rh001_049_015-    i_049    tia_h_in_001_015-    430624.8648152983
Rh001_050_015+    i_050    tia_h_in_001_015+    96468.98844157063
Rh001_050_015-    i_050    tia_h_in_001_015-    1185311.0409403413
Rh001_051_015+    i_051    tia_h_in_001_015+    853965.182210534
Rh001_051_015-    i_051    tia_h_in_001_015-    1185544.5081262991
Rh001_052_015+    i_052    tia_h_in_001_015+    349190.7130399444
Rh001_052_015-    i_052    tia_h_in_001_015-    1209270.6367251894
Rh001_053_015+    i_053    tia_h_in_001_015+    72193.78702659822
Rh001_053_015-    i_053    tia_h_in_001_015-    1203930.6840808566
Rh001_054_015+    i_054    tia_h_in_001_015+    89486.63348070974
Rh001_054_015-    i_054    tia_h_in_001_015-    1186799.3848852857
Rh001_055_015+    i_055    tia_h_in_001_015+    85141.80578483804
Rh001_055_015-    i_055    tia_h_in_001_015-    1191204.9939682214
Rh001_056_015+    i_056    tia_h_in_001_015+    1182601.7700827946
Rh001_056_015-    i_056    tia_h_in_001_015-    276668.7658803088
Rh001_057_015+    i_057    tia_h_in_001_015+    1204930.8453029727
Rh001_057_015-    i_057    tia_h_in_001_015-    726038.9667731615
Rh001_058_015+    i_058    tia_h_in_001_015+    311950.71869436087
Rh001_058_015-    i_058    tia_h_in_001_015-    1197838.2509390027
Rh001_059_015+    i_059    tia_h_in_001_015+    70321.00806203358
Rh001_059_015-    i_059    tia_h_in_001_015-    1195965.8777782505
Rh001_060_015+    i_060    tia_h_in_001_015+    131649.15635259775
Rh001_060_015-    i_060    tia_h_in_001_015-    1202984.7885245
Rh001_061_015+    i_061    tia_h_in_001_015+    1195557.0276991373
Rh001_061_015-    i_061    tia_h_in_001_015-    654773.0042948168
Rh001_062_015+    i_062    tia_h_in_001_015+    157584.74531706027
Rh001_062_015-    i_062    tia_h_in_001_015-    1205398.1343537166
Rh001_063_015+    i_063    tia_h_in_001_015+    1197374.8880320122
Rh001_063_015-    i_063    tia_h_in_001_015-    461797.82691429846
Rh001_064_015+    i_064    tia_h_in_001_015+    203115.16328553084
Rh001_064_015-    i_064    tia_h_in_001_015-    1186126.4592146522

* Neuron 16
Rh001_001_016+    i_001    tia_h_in_001_016+    32082.465029450323
Rh001_001_016-    i_001    tia_h_in_001_016-    1194984.1755900215
Rh001_002_016+    i_002    tia_h_in_001_016+    28547.81012366133
Rh001_002_016-    i_002    tia_h_in_001_016-    1203262.8948172806
Rh001_003_016+    i_003    tia_h_in_001_016+    90653.13272236873
Rh001_003_016-    i_003    tia_h_in_001_016-    1173147.9182366699
Rh001_004_016+    i_004    tia_h_in_001_016+    1178707.732457774
Rh001_004_016-    i_004    tia_h_in_001_016-    133527.81068709982
Rh001_005_016+    i_005    tia_h_in_001_016+    1197616.8987838528
Rh001_005_016-    i_005    tia_h_in_001_016-    34221.51603158376
Rh001_006_016+    i_006    tia_h_in_001_016+    1193599.6726897405
Rh001_006_016-    i_006    tia_h_in_001_016-    28801.30941548865
Rh001_007_016+    i_007    tia_h_in_001_016+    182092.44314726943
Rh001_007_016-    i_007    tia_h_in_001_016-    1194562.2491789353
Rh001_008_016+    i_008    tia_h_in_001_016+    44773.688666253176
Rh001_008_016-    i_008    tia_h_in_001_016-    1192831.1839029437
Rh001_009_016+    i_009    tia_h_in_001_016+    689702.485879857
Rh001_009_016-    i_009    tia_h_in_001_016-    1223052.154396477
Rh001_010_016+    i_010    tia_h_in_001_016+    1206671.419693078
Rh001_010_016-    i_010    tia_h_in_001_016-    204466.1586412612
Rh001_011_016+    i_011    tia_h_in_001_016+    1204248.5174702029
Rh001_011_016-    i_011    tia_h_in_001_016-    196464.48483800882
Rh001_012_016+    i_012    tia_h_in_001_016+    1206451.7139189306
Rh001_012_016-    i_012    tia_h_in_001_016-    154221.54979213982
Rh001_013_016+    i_013    tia_h_in_001_016+    237067.4167167307
Rh001_013_016-    i_013    tia_h_in_001_016-    1207494.5859171054
Rh001_014_016+    i_014    tia_h_in_001_016+    102684.95498646874
Rh001_014_016-    i_014    tia_h_in_001_016-    1195201.0892642029
Rh001_015_016+    i_015    tia_h_in_001_016+    54892.10257865244
Rh001_015_016-    i_015    tia_h_in_001_016-    1201975.9091003058
Rh001_016_016+    i_016    tia_h_in_001_016+    45318.22944119239
Rh001_016_016-    i_016    tia_h_in_001_016-    1186489.3250289597
Rh001_017_016+    i_017    tia_h_in_001_016+    164409.29558016465
Rh001_017_016-    i_017    tia_h_in_001_016-    1217988.1725956018
Rh001_018_016+    i_018    tia_h_in_001_016+    51094.40476232881
Rh001_018_016-    i_018    tia_h_in_001_016-    1198575.6134148864
Rh001_019_016+    i_019    tia_h_in_001_016+    176072.78542063234
Rh001_019_016-    i_019    tia_h_in_001_016-    1204870.1268845005
Rh001_020_016+    i_020    tia_h_in_001_016+    1193224.3855767604
Rh001_020_016-    i_020    tia_h_in_001_016-    209697.61081311078
Rh001_021_016+    i_021    tia_h_in_001_016+    1200573.8377914946
Rh001_021_016-    i_021    tia_h_in_001_016-    81668.1020677203
Rh001_022_016+    i_022    tia_h_in_001_016+    139959.78343105555
Rh001_022_016-    i_022    tia_h_in_001_016-    1188271.1964135214
Rh001_023_016+    i_023    tia_h_in_001_016+    1207776.925660858
Rh001_023_016-    i_023    tia_h_in_001_016-    894756.4300441528
Rh001_024_016+    i_024    tia_h_in_001_016+    66607.37559285211
Rh001_024_016-    i_024    tia_h_in_001_016-    1206756.3182055454
Rh001_025_016+    i_025    tia_h_in_001_016+    92175.87856791898
Rh001_025_016-    i_025    tia_h_in_001_016-    1191600.9466520152
Rh001_026_016+    i_026    tia_h_in_001_016+    1190474.0406267215
Rh001_026_016-    i_026    tia_h_in_001_016-    887838.7321871008
Rh001_027_016+    i_027    tia_h_in_001_016+    667132.5625267216
Rh001_027_016-    i_027    tia_h_in_001_016-    1191894.7326621877
Rh001_028_016+    i_028    tia_h_in_001_016+    205187.22742157005
Rh001_028_016-    i_028    tia_h_in_001_016-    1190581.644918425
Rh001_029_016+    i_029    tia_h_in_001_016+    134404.3276752817
Rh001_029_016-    i_029    tia_h_in_001_016-    1217882.93718006
Rh001_030_016+    i_030    tia_h_in_001_016+    207831.0703225506
Rh001_030_016-    i_030    tia_h_in_001_016-    1185865.1707502343
Rh001_031_016+    i_031    tia_h_in_001_016+    56728.18793565189
Rh001_031_016-    i_031    tia_h_in_001_016-    1193243.6596068763
Rh001_032_016+    i_032    tia_h_in_001_016+    65505.239009120436
Rh001_032_016-    i_032    tia_h_in_001_016-    1201378.682421145
Rh001_033_016+    i_033    tia_h_in_001_016+    132889.57874820387
Rh001_033_016-    i_033    tia_h_in_001_016-    1188400.867685365
Rh001_034_016+    i_034    tia_h_in_001_016+    127838.83031103185
Rh001_034_016-    i_034    tia_h_in_001_016-    1217889.7420553467
Rh001_035_016+    i_035    tia_h_in_001_016+    1188930.1019853777
Rh001_035_016-    i_035    tia_h_in_001_016-    148881.6042224217
Rh001_036_016+    i_036    tia_h_in_001_016+    1188319.7366166234
Rh001_036_016-    i_036    tia_h_in_001_016-    101441.92763433514
Rh001_037_016+    i_037    tia_h_in_001_016+    85268.02614745243
Rh001_037_016-    i_037    tia_h_in_001_016-    1201051.9285074829
Rh001_038_016+    i_038    tia_h_in_001_016+    42670.8867146431
Rh001_038_016-    i_038    tia_h_in_001_016-    1199217.2634933286
Rh001_039_016+    i_039    tia_h_in_001_016+    92039.32223578858
Rh001_039_016-    i_039    tia_h_in_001_016-    1194034.7354217581
Rh001_040_016+    i_040    tia_h_in_001_016+    47207.8886636882
Rh001_040_016-    i_040    tia_h_in_001_016-    1199512.107833189
Rh001_041_016+    i_041    tia_h_in_001_016+    1197884.3358004543
Rh001_041_016-    i_041    tia_h_in_001_016-    152254.30705587988
Rh001_042_016+    i_042    tia_h_in_001_016+    1198284.9494347181
Rh001_042_016-    i_042    tia_h_in_001_016-    748200.056957194
Rh001_043_016+    i_043    tia_h_in_001_016+    323902.97849930177
Rh001_043_016-    i_043    tia_h_in_001_016-    1192444.0416246897
Rh001_044_016+    i_044    tia_h_in_001_016+    45311.25158546729
Rh001_044_016-    i_044    tia_h_in_001_016-    1197468.2677980266
Rh001_045_016+    i_045    tia_h_in_001_016+    42707.56435088921
Rh001_045_016-    i_045    tia_h_in_001_016-    1195870.307074424
Rh001_046_016+    i_046    tia_h_in_001_016+    49116.12719071532
Rh001_046_016-    i_046    tia_h_in_001_016-    1194359.0687467658
Rh001_047_016+    i_047    tia_h_in_001_016+    82564.03355307919
Rh001_047_016-    i_047    tia_h_in_001_016-    1196511.1154587572
Rh001_048_016+    i_048    tia_h_in_001_016+    1196087.578424213
Rh001_048_016-    i_048    tia_h_in_001_016-    111886.81445811744
Rh001_049_016+    i_049    tia_h_in_001_016+    1206281.5932405232
Rh001_049_016-    i_049    tia_h_in_001_016-    962751.2175657691
Rh001_050_016+    i_050    tia_h_in_001_016+    1194226.2012513082
Rh001_050_016-    i_050    tia_h_in_001_016-    120114.83845264949
Rh001_051_016+    i_051    tia_h_in_001_016+    1196021.083288353
Rh001_051_016-    i_051    tia_h_in_001_016-    248847.58850301793
Rh001_052_016+    i_052    tia_h_in_001_016+    65699.74315927428
Rh001_052_016-    i_052    tia_h_in_001_016-    1206783.9492235656
Rh001_053_016+    i_053    tia_h_in_001_016+    59189.987782373435
Rh001_053_016-    i_053    tia_h_in_001_016-    1219371.8978988354
Rh001_054_016+    i_054    tia_h_in_001_016+    36441.6717634584
Rh001_054_016-    i_054    tia_h_in_001_016-    1204416.4283862354
Rh001_055_016+    i_055    tia_h_in_001_016+    61857.65615652387
Rh001_055_016-    i_055    tia_h_in_001_016-    1198351.241864108
Rh001_056_016+    i_056    tia_h_in_001_016+    1197889.2365915854
Rh001_056_016-    i_056    tia_h_in_001_016-    433256.19808061613
Rh001_057_016+    i_057    tia_h_in_001_016+    1200239.1719219699
Rh001_057_016-    i_057    tia_h_in_001_016-    129438.40776829085
Rh001_058_016+    i_058    tia_h_in_001_016+    1184439.234821575
Rh001_058_016-    i_058    tia_h_in_001_016-    1187458.8272519624
Rh001_059_016+    i_059    tia_h_in_001_016+    32284.10470018426
Rh001_059_016-    i_059    tia_h_in_001_016-    1190243.1268225554
Rh001_060_016+    i_060    tia_h_in_001_016+    26250.62502570009
Rh001_060_016-    i_060    tia_h_in_001_016-    1207907.2912045442
Rh001_061_016+    i_061    tia_h_in_001_016+    29323.262472912327
Rh001_061_016-    i_061    tia_h_in_001_016-    1210950.0589175557
Rh001_062_016+    i_062    tia_h_in_001_016+    170683.41143886573
Rh001_062_016-    i_062    tia_h_in_001_016-    1183018.8399402546
Rh001_063_016+    i_063    tia_h_in_001_016+    1200077.7934724432
Rh001_063_016-    i_063    tia_h_in_001_016-    48319.815984107736
Rh001_064_016+    i_064    tia_h_in_001_016+    1194742.0474828193
Rh001_064_016-    i_064    tia_h_in_001_016-    43305.67863537407

* Neuron 17
Rh001_001_017+    i_001    tia_h_in_001_017+    1211918.5392386662
Rh001_001_017-    i_001    tia_h_in_001_017-    178823.85218045354
Rh001_002_017+    i_002    tia_h_in_001_017+    87714.69248820175
Rh001_002_017-    i_002    tia_h_in_001_017-    1190193.1056010162
Rh001_003_017+    i_003    tia_h_in_001_017+    1198112.4019132683
Rh001_003_017-    i_003    tia_h_in_001_017-    66733.20400576602
Rh001_004_017+    i_004    tia_h_in_001_017+    1201232.9490784013
Rh001_004_017-    i_004    tia_h_in_001_017-    19885.419690492894
Rh001_005_017+    i_005    tia_h_in_001_017+    1204312.3246020824
Rh001_005_017-    i_005    tia_h_in_001_017-    104459.17109880073
Rh001_006_017+    i_006    tia_h_in_001_017+    42842.1739156243
Rh001_006_017-    i_006    tia_h_in_001_017-    1195768.1687696194
Rh001_007_017+    i_007    tia_h_in_001_017+    35905.26066118874
Rh001_007_017-    i_007    tia_h_in_001_017-    1203730.107010208
Rh001_008_017+    i_008    tia_h_in_001_017+    36061.30457836237
Rh001_008_017-    i_008    tia_h_in_001_017-    1198086.0646907918
Rh001_009_017+    i_009    tia_h_in_001_017+    418404.3050638116
Rh001_009_017-    i_009    tia_h_in_001_017-    1195303.8140754008
Rh001_010_017+    i_010    tia_h_in_001_017+    1190174.2468047764
Rh001_010_017-    i_010    tia_h_in_001_017-    131587.80918693877
Rh001_011_017+    i_011    tia_h_in_001_017+    1187295.6653756395
Rh001_011_017-    i_011    tia_h_in_001_017-    55523.47708634589
Rh001_012_017+    i_012    tia_h_in_001_017+    1183045.7637872626
Rh001_012_017-    i_012    tia_h_in_001_017-    259110.5831523522
Rh001_013_017+    i_013    tia_h_in_001_017+    61311.64708337937
Rh001_013_017-    i_013    tia_h_in_001_017-    1206188.7328577254
Rh001_014_017+    i_014    tia_h_in_001_017+    27952.76217134005
Rh001_014_017-    i_014    tia_h_in_001_017-    1202912.194641805
Rh001_015_017+    i_015    tia_h_in_001_017+    85382.46210157606
Rh001_015_017-    i_015    tia_h_in_001_017-    1193783.9864703687
Rh001_016_017+    i_016    tia_h_in_001_017+    185885.25347354813
Rh001_016_017-    i_016    tia_h_in_001_017-    1203056.6635087454
Rh001_017_017+    i_017    tia_h_in_001_017+    252852.39554609533
Rh001_017_017-    i_017    tia_h_in_001_017-    1196613.0146642926
Rh001_018_017+    i_018    tia_h_in_001_017+    1185178.12323416
Rh001_018_017-    i_018    tia_h_in_001_017-    309031.24637180095
Rh001_019_017+    i_019    tia_h_in_001_017+    1203666.0089735957
Rh001_019_017-    i_019    tia_h_in_001_017-    77917.59878829125
Rh001_020_017+    i_020    tia_h_in_001_017+    165596.41446986503
Rh001_020_017-    i_020    tia_h_in_001_017-    1212467.6654061086
Rh001_021_017+    i_021    tia_h_in_001_017+    49886.50380029054
Rh001_021_017-    i_021    tia_h_in_001_017-    1212675.9660808777
Rh001_022_017+    i_022    tia_h_in_001_017+    72423.4169820083
Rh001_022_017-    i_022    tia_h_in_001_017-    1198267.024712891
Rh001_023_017+    i_023    tia_h_in_001_017+    59381.46337950789
Rh001_023_017-    i_023    tia_h_in_001_017-    1199243.1939343137
Rh001_024_017+    i_024    tia_h_in_001_017+    1182120.4864807555
Rh001_024_017-    i_024    tia_h_in_001_017-    200345.46460503677
Rh001_025_017+    i_025    tia_h_in_001_017+    89519.49737644262
Rh001_025_017-    i_025    tia_h_in_001_017-    1185548.7154704873
Rh001_026_017+    i_026    tia_h_in_001_017+    89789.87924751395
Rh001_026_017-    i_026    tia_h_in_001_017-    1173750.5558995644
Rh001_027_017+    i_027    tia_h_in_001_017+    60340.91734850728
Rh001_027_017-    i_027    tia_h_in_001_017-    1181844.9902390644
Rh001_028_017+    i_028    tia_h_in_001_017+    36216.146657903286
Rh001_028_017-    i_028    tia_h_in_001_017-    1198405.6620979977
Rh001_029_017+    i_029    tia_h_in_001_017+    22419.821280812826
Rh001_029_017-    i_029    tia_h_in_001_017-    1208391.6498936622
Rh001_030_017+    i_030    tia_h_in_001_017+    45359.64640511235
Rh001_030_017-    i_030    tia_h_in_001_017-    1198419.3692988975
Rh001_031_017+    i_031    tia_h_in_001_017+    1193567.283479119
Rh001_031_017-    i_031    tia_h_in_001_017-    67233.4584973139
Rh001_032_017+    i_032    tia_h_in_001_017+    1213561.8383004905
Rh001_032_017-    i_032    tia_h_in_001_017-    1001685.4621879566
Rh001_033_017+    i_033    tia_h_in_001_017+    337440.07520249055
Rh001_033_017-    i_033    tia_h_in_001_017-    1217918.3805348722
Rh001_034_017+    i_034    tia_h_in_001_017+    1179674.274481998
Rh001_034_017-    i_034    tia_h_in_001_017-    52343.92740837144
Rh001_035_017+    i_035    tia_h_in_001_017+    31502.070720516793
Rh001_035_017-    i_035    tia_h_in_001_017-    1179532.871102971
Rh001_036_017+    i_036    tia_h_in_001_017+    25697.938800149986
Rh001_036_017-    i_036    tia_h_in_001_017-    1190462.8834169244
Rh001_037_017+    i_037    tia_h_in_001_017+    45534.218940575156
Rh001_037_017-    i_037    tia_h_in_001_017-    1192947.0004874861
Rh001_038_017+    i_038    tia_h_in_001_017+    83365.74385747687
Rh001_038_017-    i_038    tia_h_in_001_017-    1196692.2002278883
Rh001_039_017+    i_039    tia_h_in_001_017+    373060.4659128002
Rh001_039_017-    i_039    tia_h_in_001_017-    1206762.15739435
Rh001_040_017+    i_040    tia_h_in_001_017+    65899.60475678385
Rh001_040_017-    i_040    tia_h_in_001_017-    1178672.5605752806
Rh001_041_017+    i_041    tia_h_in_001_017+    81102.38672678523
Rh001_041_017-    i_041    tia_h_in_001_017-    1195775.028713729
Rh001_042_017+    i_042    tia_h_in_001_017+    57301.064503704874
Rh001_042_017-    i_042    tia_h_in_001_017-    1192568.0036172224
Rh001_043_017+    i_043    tia_h_in_001_017+    67851.3949074358
Rh001_043_017-    i_043    tia_h_in_001_017-    1204946.5888327507
Rh001_044_017+    i_044    tia_h_in_001_017+    78916.57739370425
Rh001_044_017-    i_044    tia_h_in_001_017-    1186754.9665445543
Rh001_045_017+    i_045    tia_h_in_001_017+    1215805.7542081259
Rh001_045_017-    i_045    tia_h_in_001_017-    549492.3588414635
Rh001_046_017+    i_046    tia_h_in_001_017+    1181188.4126946016
Rh001_046_017-    i_046    tia_h_in_001_017-    84391.70105682874
Rh001_047_017+    i_047    tia_h_in_001_017+    542041.4944061289
Rh001_047_017-    i_047    tia_h_in_001_017-    1192252.6352929797
Rh001_048_017+    i_048    tia_h_in_001_017+    156209.7000607381
Rh001_048_017-    i_048    tia_h_in_001_017-    1195196.3252689333
Rh001_049_017+    i_049    tia_h_in_001_017+    1202005.397975941
Rh001_049_017-    i_049    tia_h_in_001_017-    403053.2176312049
Rh001_050_017+    i_050    tia_h_in_001_017+    75753.27859935412
Rh001_050_017-    i_050    tia_h_in_001_017-    1198647.3972957784
Rh001_051_017+    i_051    tia_h_in_001_017+    47922.589535265404
Rh001_051_017-    i_051    tia_h_in_001_017-    1206917.1214361333
Rh001_052_017+    i_052    tia_h_in_001_017+    53082.59019923191
Rh001_052_017-    i_052    tia_h_in_001_017-    1179998.2967931004
Rh001_053_017+    i_053    tia_h_in_001_017+    553172.759853237
Rh001_053_017-    i_053    tia_h_in_001_017-    1192885.7584912635
Rh001_054_017+    i_054    tia_h_in_001_017+    1195002.3335362026
Rh001_054_017-    i_054    tia_h_in_001_017-    50275.044033199774
Rh001_055_017+    i_055    tia_h_in_001_017+    1200091.0526604573
Rh001_055_017-    i_055    tia_h_in_001_017-    263544.0463735307
Rh001_056_017+    i_056    tia_h_in_001_017+    1203839.363050108
Rh001_056_017-    i_056    tia_h_in_001_017-    107521.0337869835
Rh001_057_017+    i_057    tia_h_in_001_017+    48018.35383722754
Rh001_057_017-    i_057    tia_h_in_001_017-    1222318.8745592528
Rh001_058_017+    i_058    tia_h_in_001_017+    37436.46413755729
Rh001_058_017-    i_058    tia_h_in_001_017-    1191599.6856686817
Rh001_059_017+    i_059    tia_h_in_001_017+    42121.14829177433
Rh001_059_017-    i_059    tia_h_in_001_017-    1201884.6702618639
Rh001_060_017+    i_060    tia_h_in_001_017+    1214765.8396998756
Rh001_060_017-    i_060    tia_h_in_001_017-    72132.78393716048
Rh001_061_017+    i_061    tia_h_in_001_017+    1218684.560834335
Rh001_061_017-    i_061    tia_h_in_001_017-    21297.475575343815
Rh001_062_017+    i_062    tia_h_in_001_017+    1193747.0683608055
Rh001_062_017-    i_062    tia_h_in_001_017-    73558.73664458847
Rh001_063_017+    i_063    tia_h_in_001_017+    65585.54074947884
Rh001_063_017-    i_063    tia_h_in_001_017-    1196364.6506853155
Rh001_064_017+    i_064    tia_h_in_001_017+    116736.92585225144
Rh001_064_017-    i_064    tia_h_in_001_017-    1201723.1321462

* Neuron 18
Rh001_001_018+    i_001    tia_h_in_001_018+    1194931.5455403586
Rh001_001_018-    i_001    tia_h_in_001_018-    64473.307036160055
Rh001_002_018+    i_002    tia_h_in_001_018+    1201772.5599831217
Rh001_002_018-    i_002    tia_h_in_001_018-    58353.840783387
Rh001_003_018+    i_003    tia_h_in_001_018+    331860.0012895194
Rh001_003_018-    i_003    tia_h_in_001_018-    1187893.0778214794
Rh001_004_018+    i_004    tia_h_in_001_018+    1211608.7622008303
Rh001_004_018-    i_004    tia_h_in_001_018-    629040.3561755971
Rh001_005_018+    i_005    tia_h_in_001_018+    135436.0991526353
Rh001_005_018-    i_005    tia_h_in_001_018-    1198496.4547014907
Rh001_006_018+    i_006    tia_h_in_001_018+    1201099.0619992614
Rh001_006_018-    i_006    tia_h_in_001_018-    949903.084844214
Rh001_007_018+    i_007    tia_h_in_001_018+    95486.07411985353
Rh001_007_018-    i_007    tia_h_in_001_018-    1208762.6489867026
Rh001_008_018+    i_008    tia_h_in_001_018+    63251.80171387023
Rh001_008_018-    i_008    tia_h_in_001_018-    1207523.4051983624
Rh001_009_018+    i_009    tia_h_in_001_018+    1205610.9971962466
Rh001_009_018-    i_009    tia_h_in_001_018-    97129.12746100349
Rh001_010_018+    i_010    tia_h_in_001_018+    1206651.498874643
Rh001_010_018-    i_010    tia_h_in_001_018-    593758.5858684505
Rh001_011_018+    i_011    tia_h_in_001_018+    70909.87183720001
Rh001_011_018-    i_011    tia_h_in_001_018-    1198792.5273510488
Rh001_012_018+    i_012    tia_h_in_001_018+    70527.87303838399
Rh001_012_018-    i_012    tia_h_in_001_018-    1197015.2762698263
Rh001_013_018+    i_013    tia_h_in_001_018+    153059.01202137003
Rh001_013_018-    i_013    tia_h_in_001_018-    1185105.099714851
Rh001_014_018+    i_014    tia_h_in_001_018+    66975.41013117299
Rh001_014_018-    i_014    tia_h_in_001_018-    1199673.109750015
Rh001_015_018+    i_015    tia_h_in_001_018+    77793.6240778753
Rh001_015_018-    i_015    tia_h_in_001_018-    1206463.697077086
Rh001_016_018+    i_016    tia_h_in_001_018+    1181166.147651845
Rh001_016_018-    i_016    tia_h_in_001_018-    190012.37201954078
Rh001_017_018+    i_017    tia_h_in_001_018+    101830.0480464846
Rh001_017_018-    i_017    tia_h_in_001_018-    1200974.1568312463
Rh001_018_018+    i_018    tia_h_in_001_018+    82043.81434589004
Rh001_018_018-    i_018    tia_h_in_001_018-    1193528.0369691907
Rh001_019_018+    i_019    tia_h_in_001_018+    68667.15434816596
Rh001_019_018-    i_019    tia_h_in_001_018-    1215198.4113685759
Rh001_020_018+    i_020    tia_h_in_001_018+    1192340.483304392
Rh001_020_018-    i_020    tia_h_in_001_018-    989757.2184263339
Rh001_021_018+    i_021    tia_h_in_001_018+    91216.46521964739
Rh001_021_018-    i_021    tia_h_in_001_018-    1211713.4424882666
Rh001_022_018+    i_022    tia_h_in_001_018+    157737.79575379076
Rh001_022_018-    i_022    tia_h_in_001_018-    1200478.2479816352
Rh001_023_018+    i_023    tia_h_in_001_018+    226381.37167262982
Rh001_023_018-    i_023    tia_h_in_001_018-    1201256.5446171209
Rh001_024_018+    i_024    tia_h_in_001_018+    118022.89163581711
Rh001_024_018-    i_024    tia_h_in_001_018-    1193028.4739294203
Rh001_025_018+    i_025    tia_h_in_001_018+    75051.87069582936
Rh001_025_018-    i_025    tia_h_in_001_018-    1196471.4453431095
Rh001_026_018+    i_026    tia_h_in_001_018+    51291.53682543977
Rh001_026_018-    i_026    tia_h_in_001_018-    1195241.372923051
Rh001_027_018+    i_027    tia_h_in_001_018+    68818.75257913917
Rh001_027_018-    i_027    tia_h_in_001_018-    1208465.283518185
Rh001_028_018+    i_028    tia_h_in_001_018+    61743.83650655765
Rh001_028_018-    i_028    tia_h_in_001_018-    1185543.809060514
Rh001_029_018+    i_029    tia_h_in_001_018+    1189902.938501206
Rh001_029_018-    i_029    tia_h_in_001_018-    206746.238452938
Rh001_030_018+    i_030    tia_h_in_001_018+    1201448.6244971787
Rh001_030_018-    i_030    tia_h_in_001_018-    162274.44206656338
Rh001_031_018+    i_031    tia_h_in_001_018+    51880.56134674794
Rh001_031_018-    i_031    tia_h_in_001_018-    1209098.8621849888
Rh001_032_018+    i_032    tia_h_in_001_018+    183739.56509448035
Rh001_032_018-    i_032    tia_h_in_001_018-    1219398.5816731935
Rh001_033_018+    i_033    tia_h_in_001_018+    41090.434350770774
Rh001_033_018-    i_033    tia_h_in_001_018-    1193270.910609933
Rh001_034_018+    i_034    tia_h_in_001_018+    60899.62066168207
Rh001_034_018-    i_034    tia_h_in_001_018-    1205108.9254370152
Rh001_035_018+    i_035    tia_h_in_001_018+    251610.64041755756
Rh001_035_018-    i_035    tia_h_in_001_018-    1205453.5661352065
Rh001_036_018+    i_036    tia_h_in_001_018+    76192.49020627145
Rh001_036_018-    i_036    tia_h_in_001_018-    1191633.1959728557
Rh001_037_018+    i_037    tia_h_in_001_018+    66347.25787250968
Rh001_037_018-    i_037    tia_h_in_001_018-    1189358.1150544505
Rh001_038_018+    i_038    tia_h_in_001_018+    55794.15829111854
Rh001_038_018-    i_038    tia_h_in_001_018-    1204916.8300659305
Rh001_039_018+    i_039    tia_h_in_001_018+    71529.65863581195
Rh001_039_018-    i_039    tia_h_in_001_018-    1199568.8229650212
Rh001_040_018+    i_040    tia_h_in_001_018+    26921.54768007599
Rh001_040_018-    i_040    tia_h_in_001_018-    1201962.8008240946
Rh001_041_018+    i_041    tia_h_in_001_018+    283123.35995278554
Rh001_041_018-    i_041    tia_h_in_001_018-    1197211.2946625238
Rh001_042_018+    i_042    tia_h_in_001_018+    1169831.863722146
Rh001_042_018-    i_042    tia_h_in_001_018-    1191509.457810939
Rh001_043_018+    i_043    tia_h_in_001_018+    165017.64820708949
Rh001_043_018-    i_043    tia_h_in_001_018-    1190386.8635157545
Rh001_044_018+    i_044    tia_h_in_001_018+    139623.23911613945
Rh001_044_018-    i_044    tia_h_in_001_018-    1186162.023371547
Rh001_045_018+    i_045    tia_h_in_001_018+    234037.5010844867
Rh001_045_018-    i_045    tia_h_in_001_018-    1205291.2924606265
Rh001_046_018+    i_046    tia_h_in_001_018+    40455.46228190769
Rh001_046_018-    i_046    tia_h_in_001_018-    1180518.136259158
Rh001_047_018+    i_047    tia_h_in_001_018+    51692.515682157646
Rh001_047_018-    i_047    tia_h_in_001_018-    1197271.42293977
Rh001_048_018+    i_048    tia_h_in_001_018+    41857.1945583611
Rh001_048_018-    i_048    tia_h_in_001_018-    1204593.5822199953
Rh001_049_018+    i_049    tia_h_in_001_018+    195516.62141558094
Rh001_049_018-    i_049    tia_h_in_001_018-    1204562.541927114
Rh001_050_018+    i_050    tia_h_in_001_018+    112910.18752358195
Rh001_050_018-    i_050    tia_h_in_001_018-    1211102.491779387
Rh001_051_018+    i_051    tia_h_in_001_018+    289632.35063015914
Rh001_051_018-    i_051    tia_h_in_001_018-    1198653.7897138165
Rh001_052_018+    i_052    tia_h_in_001_018+    420005.3921557324
Rh001_052_018-    i_052    tia_h_in_001_018-    1200802.937810007
Rh001_053_018+    i_053    tia_h_in_001_018+    197709.49188560317
Rh001_053_018-    i_053    tia_h_in_001_018-    1201655.3498302521
Rh001_054_018+    i_054    tia_h_in_001_018+    1025847.1066129416
Rh001_054_018-    i_054    tia_h_in_001_018-    1191372.5023374488
Rh001_055_018+    i_055    tia_h_in_001_018+    81644.48028613583
Rh001_055_018-    i_055    tia_h_in_001_018-    1198687.222822294
Rh001_056_018+    i_056    tia_h_in_001_018+    1186818.91403566
Rh001_056_018-    i_056    tia_h_in_001_018-    36968.98124732966
Rh001_057_018+    i_057    tia_h_in_001_018+    77977.98916936362
Rh001_057_018-    i_057    tia_h_in_001_018-    1199091.5247024428
Rh001_058_018+    i_058    tia_h_in_001_018+    106913.14303110639
Rh001_058_018-    i_058    tia_h_in_001_018-    1197759.2340232797
Rh001_059_018+    i_059    tia_h_in_001_018+    375564.8468822015
Rh001_059_018-    i_059    tia_h_in_001_018-    1190434.8306590142
Rh001_060_018+    i_060    tia_h_in_001_018+    52203.8600134831
Rh001_060_018-    i_060    tia_h_in_001_018-    1187217.1948122692
Rh001_061_018+    i_061    tia_h_in_001_018+    343347.56143649865
Rh001_061_018-    i_061    tia_h_in_001_018-    1191293.7580021424
Rh001_062_018+    i_062    tia_h_in_001_018+    1220636.6458233253
Rh001_062_018-    i_062    tia_h_in_001_018-    186768.80638673782
Rh001_063_018+    i_063    tia_h_in_001_018+    1206517.633466925
Rh001_063_018-    i_063    tia_h_in_001_018-    26871.064110130912
Rh001_064_018+    i_064    tia_h_in_001_018+    1186901.4949452274
Rh001_064_018-    i_064    tia_h_in_001_018-    46490.85600339946

* Neuron 19
Rh001_001_019+    i_001    tia_h_in_001_019+    55739.49102623571
Rh001_001_019-    i_001    tia_h_in_001_019-    1224528.9436101778
Rh001_002_019+    i_002    tia_h_in_001_019+    56612.45808353101
Rh001_002_019-    i_002    tia_h_in_001_019-    1213655.638142121
Rh001_003_019+    i_003    tia_h_in_001_019+    24102.58466290939
Rh001_003_019-    i_003    tia_h_in_001_019-    1203695.2679412623
Rh001_004_019+    i_004    tia_h_in_001_019+    90782.63934471317
Rh001_004_019-    i_004    tia_h_in_001_019-    1205443.9344062975
Rh001_005_019+    i_005    tia_h_in_001_019+    1196197.8747179534
Rh001_005_019-    i_005    tia_h_in_001_019-    111613.77332760674
Rh001_006_019+    i_006    tia_h_in_001_019+    1197347.6587093228
Rh001_006_019-    i_006    tia_h_in_001_019-    62850.6844809924
Rh001_007_019+    i_007    tia_h_in_001_019+    1207359.0777138073
Rh001_007_019-    i_007    tia_h_in_001_019-    238476.2090894461
Rh001_008_019+    i_008    tia_h_in_001_019+    1215992.3913811739
Rh001_008_019-    i_008    tia_h_in_001_019-    111855.05661816007
Rh001_009_019+    i_009    tia_h_in_001_019+    79750.93969363098
Rh001_009_019-    i_009    tia_h_in_001_019-    1207645.2092339194
Rh001_010_019+    i_010    tia_h_in_001_019+    44512.50296485872
Rh001_010_019-    i_010    tia_h_in_001_019-    1192067.1525362697
Rh001_011_019+    i_011    tia_h_in_001_019+    443703.7991495319
Rh001_011_019-    i_011    tia_h_in_001_019-    1193619.4616741173
Rh001_012_019+    i_012    tia_h_in_001_019+    1210001.2959793978
Rh001_012_019-    i_012    tia_h_in_001_019-    89335.13179574534
Rh001_013_019+    i_013    tia_h_in_001_019+    1190892.863276322
Rh001_013_019-    i_013    tia_h_in_001_019-    177396.66995117083
Rh001_014_019+    i_014    tia_h_in_001_019+    322644.43889498495
Rh001_014_019-    i_014    tia_h_in_001_019-    1215386.7982567782
Rh001_015_019+    i_015    tia_h_in_001_019+    679440.4508944533
Rh001_015_019-    i_015    tia_h_in_001_019-    1207105.095403654
Rh001_016_019+    i_016    tia_h_in_001_019+    77921.23751845834
Rh001_016_019-    i_016    tia_h_in_001_019-    1205568.0052130008
Rh001_017_019+    i_017    tia_h_in_001_019+    37025.26185193297
Rh001_017_019-    i_017    tia_h_in_001_019-    1201747.9102017828
Rh001_018_019+    i_018    tia_h_in_001_019+    38048.97363188566
Rh001_018_019-    i_018    tia_h_in_001_019-    1194797.4758783206
Rh001_019_019+    i_019    tia_h_in_001_019+    97597.57691653025
Rh001_019_019-    i_019    tia_h_in_001_019-    1198624.7624892169
Rh001_020_019+    i_020    tia_h_in_001_019+    116633.94384500127
Rh001_020_019-    i_020    tia_h_in_001_019-    1215466.0848703382
Rh001_021_019+    i_021    tia_h_in_001_019+    1198245.5805229964
Rh001_021_019-    i_021    tia_h_in_001_019-    388123.3801699234
Rh001_022_019+    i_022    tia_h_in_001_019+    530522.4050185971
Rh001_022_019-    i_022    tia_h_in_001_019-    1206186.0181976305
Rh001_023_019+    i_023    tia_h_in_001_019+    117295.78531794834
Rh001_023_019-    i_023    tia_h_in_001_019-    1197739.5688221464
Rh001_024_019+    i_024    tia_h_in_001_019+    80995.1445931053
Rh001_024_019-    i_024    tia_h_in_001_019-    1190505.502611069
Rh001_025_019+    i_025    tia_h_in_001_019+    41348.57900741873
Rh001_025_019-    i_025    tia_h_in_001_019-    1192424.5476779619
Rh001_026_019+    i_026    tia_h_in_001_019+    103282.36023116035
Rh001_026_019-    i_026    tia_h_in_001_019-    1214099.5863884117
Rh001_027_019+    i_027    tia_h_in_001_019+    1203548.0603144749
Rh001_027_019-    i_027    tia_h_in_001_019-    205341.17996779023
Rh001_028_019+    i_028    tia_h_in_001_019+    272724.1524668868
Rh001_028_019-    i_028    tia_h_in_001_019-    1206589.3132128662
Rh001_029_019+    i_029    tia_h_in_001_019+    1221820.9835483548
Rh001_029_019-    i_029    tia_h_in_001_019-    264858.44031361304
Rh001_030_019+    i_030    tia_h_in_001_019+    1193851.8182583407
Rh001_030_019-    i_030    tia_h_in_001_019-    235002.94593389778
Rh001_031_019+    i_031    tia_h_in_001_019+    71243.1224687886
Rh001_031_019-    i_031    tia_h_in_001_019-    1204977.393297857
Rh001_032_019+    i_032    tia_h_in_001_019+    64844.18385077241
Rh001_032_019-    i_032    tia_h_in_001_019-    1202879.1419313254
Rh001_033_019+    i_033    tia_h_in_001_019+    74509.32498070036
Rh001_033_019-    i_033    tia_h_in_001_019-    1204149.428872777
Rh001_034_019+    i_034    tia_h_in_001_019+    94646.29275699386
Rh001_034_019-    i_034    tia_h_in_001_019-    1180019.7732697865
Rh001_035_019+    i_035    tia_h_in_001_019+    1195285.575396283
Rh001_035_019-    i_035    tia_h_in_001_019-    913091.4744738806
Rh001_036_019+    i_036    tia_h_in_001_019+    1176050.9442367926
Rh001_036_019-    i_036    tia_h_in_001_019-    354676.36439934286
Rh001_037_019+    i_037    tia_h_in_001_019+    1207170.5467022145
Rh001_037_019-    i_037    tia_h_in_001_019-    165310.90985120228
Rh001_038_019+    i_038    tia_h_in_001_019+    75002.10902203502
Rh001_038_019-    i_038    tia_h_in_001_019-    1185113.2017444975
Rh001_039_019+    i_039    tia_h_in_001_019+    141057.91216182543
Rh001_039_019-    i_039    tia_h_in_001_019-    1210318.1456948558
Rh001_040_019+    i_040    tia_h_in_001_019+    50889.82057567572
Rh001_040_019-    i_040    tia_h_in_001_019-    1198820.7494479981
Rh001_041_019+    i_041    tia_h_in_001_019+    1193892.4512110557
Rh001_041_019-    i_041    tia_h_in_001_019-    339199.90556540195
Rh001_042_019+    i_042    tia_h_in_001_019+    1210488.7578634822
Rh001_042_019-    i_042    tia_h_in_001_019-    387183.6224144079
Rh001_043_019+    i_043    tia_h_in_001_019+    1180585.4817226867
Rh001_043_019-    i_043    tia_h_in_001_019-    155367.9386874508
Rh001_044_019+    i_044    tia_h_in_001_019+    138852.0017262874
Rh001_044_019-    i_044    tia_h_in_001_019-    1179244.8284429787
Rh001_045_019+    i_045    tia_h_in_001_019+    70042.06737875356
Rh001_045_019-    i_045    tia_h_in_001_019-    1211804.3587281094
Rh001_046_019+    i_046    tia_h_in_001_019+    41255.18132294525
Rh001_046_019-    i_046    tia_h_in_001_019-    1216465.043861278
Rh001_047_019+    i_047    tia_h_in_001_019+    74550.16389837243
Rh001_047_019-    i_047    tia_h_in_001_019-    1207737.1295854494
Rh001_048_019+    i_048    tia_h_in_001_019+    78043.71546794788
Rh001_048_019-    i_048    tia_h_in_001_019-    1192060.182595605
Rh001_049_019+    i_049    tia_h_in_001_019+    1211230.5067858344
Rh001_049_019-    i_049    tia_h_in_001_019-    276455.12650071067
Rh001_050_019+    i_050    tia_h_in_001_019+    1209007.5211239138
Rh001_050_019-    i_050    tia_h_in_001_019-    132896.4846037451
Rh001_051_019+    i_051    tia_h_in_001_019+    1201959.0412933505
Rh001_051_019-    i_051    tia_h_in_001_019-    133829.98947677857
Rh001_052_019+    i_052    tia_h_in_001_019+    130524.4047377884
Rh001_052_019-    i_052    tia_h_in_001_019-    1198362.647226264
Rh001_053_019+    i_053    tia_h_in_001_019+    143786.81216925298
Rh001_053_019-    i_053    tia_h_in_001_019-    1202333.2959166295
Rh001_054_019+    i_054    tia_h_in_001_019+    49137.42076661252
Rh001_054_019-    i_054    tia_h_in_001_019-    1196314.847949076
Rh001_055_019+    i_055    tia_h_in_001_019+    37657.944033004314
Rh001_055_019-    i_055    tia_h_in_001_019-    1201635.5949807288
Rh001_056_019+    i_056    tia_h_in_001_019+    134272.62582467066
Rh001_056_019-    i_056    tia_h_in_001_019-    1193677.3078167513
Rh001_057_019+    i_057    tia_h_in_001_019+    1209520.4996611555
Rh001_057_019-    i_057    tia_h_in_001_019-    36218.694117381754
Rh001_058_019+    i_058    tia_h_in_001_019+    1198651.691605446
Rh001_058_019-    i_058    tia_h_in_001_019-    127205.5312955244
Rh001_059_019+    i_059    tia_h_in_001_019+    201187.20994345922
Rh001_059_019-    i_059    tia_h_in_001_019-    1195943.1614101233
Rh001_060_019+    i_060    tia_h_in_001_019+    30587.919629062766
Rh001_060_019-    i_060    tia_h_in_001_019-    1210662.4362463155
Rh001_061_019+    i_061    tia_h_in_001_019+    19979.78950102966
Rh001_061_019-    i_061    tia_h_in_001_019-    1187639.5235779828
Rh001_062_019+    i_062    tia_h_in_001_019+    35048.049529062366
Rh001_062_019-    i_062    tia_h_in_001_019-    1188150.0613397676
Rh001_063_019+    i_063    tia_h_in_001_019+    1199239.0084783833
Rh001_063_019-    i_063    tia_h_in_001_019-    252001.6408987868
Rh001_064_019+    i_064    tia_h_in_001_019+    814400.5386346555
Rh001_064_019-    i_064    tia_h_in_001_019-    1194865.325425035

* Neuron 20
Rh001_001_020+    i_001    tia_h_in_001_020+    1205329.5144089663
Rh001_001_020-    i_001    tia_h_in_001_020-    166474.33475806325
Rh001_002_020+    i_002    tia_h_in_001_020+    1186190.741968753
Rh001_002_020-    i_002    tia_h_in_001_020-    115413.20178486725
Rh001_003_020+    i_003    tia_h_in_001_020+    1197477.004299363
Rh001_003_020-    i_003    tia_h_in_001_020-    76593.38438763413
Rh001_004_020+    i_004    tia_h_in_001_020+    88911.5896736486
Rh001_004_020-    i_004    tia_h_in_001_020-    1198260.1537894618
Rh001_005_020+    i_005    tia_h_in_001_020+    151776.62525026494
Rh001_005_020-    i_005    tia_h_in_001_020-    1207181.6365442297
Rh001_006_020+    i_006    tia_h_in_001_020+    69441.11729217877
Rh001_006_020-    i_006    tia_h_in_001_020-    1202097.052487548
Rh001_007_020+    i_007    tia_h_in_001_020+    46345.16738310396
Rh001_007_020-    i_007    tia_h_in_001_020-    1185348.4092441967
Rh001_008_020+    i_008    tia_h_in_001_020+    47976.08589678611
Rh001_008_020-    i_008    tia_h_in_001_020-    1201286.2171322757
Rh001_009_020+    i_009    tia_h_in_001_020+    127143.11052423462
Rh001_009_020-    i_009    tia_h_in_001_020-    1187589.3364570362
Rh001_010_020+    i_010    tia_h_in_001_020+    1198771.571957112
Rh001_010_020-    i_010    tia_h_in_001_020-    45813.960723275195
Rh001_011_020+    i_011    tia_h_in_001_020+    36603.66894362987
Rh001_011_020-    i_011    tia_h_in_001_020-    1198226.1619526548
Rh001_012_020+    i_012    tia_h_in_001_020+    47021.81988490256
Rh001_012_020-    i_012    tia_h_in_001_020-    1196712.037851958
Rh001_013_020+    i_013    tia_h_in_001_020+    218860.6012280039
Rh001_013_020-    i_013    tia_h_in_001_020-    1191625.3901639513
Rh001_014_020+    i_014    tia_h_in_001_020+    45938.09771194488
Rh001_014_020-    i_014    tia_h_in_001_020-    1193221.5025872185
Rh001_015_020+    i_015    tia_h_in_001_020+    90309.63945345579
Rh001_015_020-    i_015    tia_h_in_001_020-    1203623.301087055
Rh001_016_020+    i_016    tia_h_in_001_020+    78267.67217727141
Rh001_016_020-    i_016    tia_h_in_001_020-    1216478.6779439729
Rh001_017_020+    i_017    tia_h_in_001_020+    1188063.8431092293
Rh001_017_020-    i_017    tia_h_in_001_020-    75582.11829330279
Rh001_018_020+    i_018    tia_h_in_001_020+    86474.11801315742
Rh001_018_020-    i_018    tia_h_in_001_020-    1211636.8958493902
Rh001_019_020+    i_019    tia_h_in_001_020+    71220.300484703
Rh001_019_020-    i_019    tia_h_in_001_020-    1185501.7339976018
Rh001_020_020+    i_020    tia_h_in_001_020+    64599.1613488992
Rh001_020_020-    i_020    tia_h_in_001_020-    1191401.2822910794
Rh001_021_020+    i_021    tia_h_in_001_020+    199413.81195423557
Rh001_021_020-    i_021    tia_h_in_001_020-    1195022.4923020538
Rh001_022_020+    i_022    tia_h_in_001_020+    211274.0863272718
Rh001_022_020-    i_022    tia_h_in_001_020-    1207048.3992028367
Rh001_023_020+    i_023    tia_h_in_001_020+    96685.547738607
Rh001_023_020-    i_023    tia_h_in_001_020-    1189070.6809804346
Rh001_024_020+    i_024    tia_h_in_001_020+    48828.98156728301
Rh001_024_020-    i_024    tia_h_in_001_020-    1209470.3087932793
Rh001_025_020+    i_025    tia_h_in_001_020+    123424.7519268589
Rh001_025_020-    i_025    tia_h_in_001_020-    1201422.3421447482
Rh001_026_020+    i_026    tia_h_in_001_020+    108575.4239869821
Rh001_026_020-    i_026    tia_h_in_001_020-    1186144.7084330602
Rh001_027_020+    i_027    tia_h_in_001_020+    321137.32687991066
Rh001_027_020-    i_027    tia_h_in_001_020-    1190891.8001729643
Rh001_028_020+    i_028    tia_h_in_001_020+    1198220.3190175146
Rh001_028_020-    i_028    tia_h_in_001_020-    89223.40432455478
Rh001_029_020+    i_029    tia_h_in_001_020+    1202011.6076494588
Rh001_029_020-    i_029    tia_h_in_001_020-    267294.17247239524
Rh001_030_020+    i_030    tia_h_in_001_020+    647553.8284474388
Rh001_030_020-    i_030    tia_h_in_001_020-    1209882.2273128196
Rh001_031_020+    i_031    tia_h_in_001_020+    1200914.4452605557
Rh001_031_020-    i_031    tia_h_in_001_020-    1079081.0479227358
Rh001_032_020+    i_032    tia_h_in_001_020+    122151.93464505886
Rh001_032_020-    i_032    tia_h_in_001_020-    1201710.0755126318
Rh001_033_020+    i_033    tia_h_in_001_020+    102624.06253261755
Rh001_033_020-    i_033    tia_h_in_001_020-    1200173.4705674993
Rh001_034_020+    i_034    tia_h_in_001_020+    237426.57220130638
Rh001_034_020-    i_034    tia_h_in_001_020-    1209280.3382480943
Rh001_035_020+    i_035    tia_h_in_001_020+    85301.46556611305
Rh001_035_020-    i_035    tia_h_in_001_020-    1201503.5909069437
Rh001_036_020+    i_036    tia_h_in_001_020+    853728.2062842617
Rh001_036_020-    i_036    tia_h_in_001_020-    1200648.157171731
Rh001_037_020+    i_037    tia_h_in_001_020+    1214933.3287877054
Rh001_037_020-    i_037    tia_h_in_001_020-    181600.2293339225
Rh001_038_020+    i_038    tia_h_in_001_020+    92567.64555410173
Rh001_038_020-    i_038    tia_h_in_001_020-    1188446.2612785446
Rh001_039_020+    i_039    tia_h_in_001_020+    78031.52778270388
Rh001_039_020-    i_039    tia_h_in_001_020-    1205402.6357238183
Rh001_040_020+    i_040    tia_h_in_001_020+    1198073.9660148714
Rh001_040_020-    i_040    tia_h_in_001_020-    248289.34433361204
Rh001_041_020+    i_041    tia_h_in_001_020+    107633.88611934143
Rh001_041_020-    i_041    tia_h_in_001_020-    1217399.734366432
Rh001_042_020+    i_042    tia_h_in_001_020+    61502.050022922806
Rh001_042_020-    i_042    tia_h_in_001_020-    1201752.3027479001
Rh001_043_020+    i_043    tia_h_in_001_020+    1174943.3772372412
Rh001_043_020-    i_043    tia_h_in_001_020-    97554.20249284092
Rh001_044_020+    i_044    tia_h_in_001_020+    1192509.490578749
Rh001_044_020-    i_044    tia_h_in_001_020-    194687.55443779714
Rh001_045_020+    i_045    tia_h_in_001_020+    92380.24294322025
Rh001_045_020-    i_045    tia_h_in_001_020-    1184114.4758908183
Rh001_046_020+    i_046    tia_h_in_001_020+    59567.1103108158
Rh001_046_020-    i_046    tia_h_in_001_020-    1203770.069284271
Rh001_047_020+    i_047    tia_h_in_001_020+    61791.107274365706
Rh001_047_020-    i_047    tia_h_in_001_020-    1207479.6870393045
Rh001_048_020+    i_048    tia_h_in_001_020+    158598.1647659511
Rh001_048_020-    i_048    tia_h_in_001_020-    1201737.7440060189
Rh001_049_020+    i_049    tia_h_in_001_020+    59613.8879454804
Rh001_049_020-    i_049    tia_h_in_001_020-    1191919.6671312724
Rh001_050_020+    i_050    tia_h_in_001_020+    108996.66742840954
Rh001_050_020-    i_050    tia_h_in_001_020-    1202075.1877760098
Rh001_051_020+    i_051    tia_h_in_001_020+    46996.42540307881
Rh001_051_020-    i_051    tia_h_in_001_020-    1195565.4676346183
Rh001_052_020+    i_052    tia_h_in_001_020+    65820.57750320484
Rh001_052_020-    i_052    tia_h_in_001_020-    1198782.678128582
Rh001_053_020+    i_053    tia_h_in_001_020+    106248.42840612023
Rh001_053_020-    i_053    tia_h_in_001_020-    1211471.4023218986
Rh001_054_020+    i_054    tia_h_in_001_020+    63604.365607066466
Rh001_054_020-    i_054    tia_h_in_001_020-    1208348.2168410057
Rh001_055_020+    i_055    tia_h_in_001_020+    1192746.7362056065
Rh001_055_020-    i_055    tia_h_in_001_020-    66845.5810352792
Rh001_056_020+    i_056    tia_h_in_001_020+    302929.2382994135
Rh001_056_020-    i_056    tia_h_in_001_020-    1215030.880705949
Rh001_057_020+    i_057    tia_h_in_001_020+    51942.36632616385
Rh001_057_020-    i_057    tia_h_in_001_020-    1211785.081485598
Rh001_058_020+    i_058    tia_h_in_001_020+    73450.4251502012
Rh001_058_020-    i_058    tia_h_in_001_020-    1199115.2246671803
Rh001_059_020+    i_059    tia_h_in_001_020+    43090.39566112174
Rh001_059_020-    i_059    tia_h_in_001_020-    1213375.313269603
Rh001_060_020+    i_060    tia_h_in_001_020+    113083.96431944132
Rh001_060_020-    i_060    tia_h_in_001_020-    1202195.2509838266
Rh001_061_020+    i_061    tia_h_in_001_020+    129374.12933397295
Rh001_061_020-    i_061    tia_h_in_001_020-    1210833.8393955126
Rh001_062_020+    i_062    tia_h_in_001_020+    1196579.438113417
Rh001_062_020-    i_062    tia_h_in_001_020-    90790.71269091305
Rh001_063_020+    i_063    tia_h_in_001_020+    1195205.8695021046
Rh001_063_020-    i_063    tia_h_in_001_020-    50785.664739993386
Rh001_064_020+    i_064    tia_h_in_001_020+    1198557.714385242
Rh001_064_020-    i_064    tia_h_in_001_020-    60018.32209251613

* ----- Bias
    
        
Rb_h001_001+    b_001    tia_h_in_001_001+    1188345.622481674
Rb_h001_001-    b_001    tia_h_in_001_001-    95922.6017438917
Rb_h001_002+    b_001    tia_h_in_001_002+    131968.6630804123
Rb_h001_002-    b_001    tia_h_in_001_002-    1198218.3393353785
Rb_h001_003+    b_001    tia_h_in_001_003+    1202015.402830119
Rb_h001_003-    b_001    tia_h_in_001_003-    68008.88550068667
Rb_h001_004+    b_001    tia_h_in_001_004+    1205139.9824855065
Rb_h001_004-    b_001    tia_h_in_001_004-    290788.22777819267
Rb_h001_005+    b_001    tia_h_in_001_005+    288058.4632485629
Rb_h001_005-    b_001    tia_h_in_001_005-    1194362.9302600855
Rb_h001_006+    b_001    tia_h_in_001_006+    566329.8875897297
Rb_h001_006-    b_001    tia_h_in_001_006-    1193029.7667044236
Rb_h001_007+    b_001    tia_h_in_001_007+    245570.174356554
Rb_h001_007-    b_001    tia_h_in_001_007-    1188360.5921319455
Rb_h001_008+    b_001    tia_h_in_001_008+    222468.67001479203
Rb_h001_008-    b_001    tia_h_in_001_008-    1192714.7333271494
Rb_h001_009+    b_001    tia_h_in_001_009+    148097.02323453352
Rb_h001_009-    b_001    tia_h_in_001_009-    1195475.3508322441
Rb_h001_010+    b_001    tia_h_in_001_010+    1205163.72196999
Rb_h001_010-    b_001    tia_h_in_001_010-    551472.7898237195
Rb_h001_011+    b_001    tia_h_in_001_011+    174161.2468905211
Rb_h001_011-    b_001    tia_h_in_001_011-    1180755.0096856372
Rb_h001_012+    b_001    tia_h_in_001_012+    120084.42003991439
Rb_h001_012-    b_001    tia_h_in_001_012-    1196864.3645694721
Rb_h001_013+    b_001    tia_h_in_001_013+    348324.3478796827
Rb_h001_013-    b_001    tia_h_in_001_013-    1213934.2054178682
Rb_h001_014+    b_001    tia_h_in_001_014+    1206364.811667164
Rb_h001_014-    b_001    tia_h_in_001_014-    291094.0596806918
Rb_h001_015+    b_001    tia_h_in_001_015+    906590.1403948745
Rb_h001_015-    b_001    tia_h_in_001_015-    1214333.4354772524
Rb_h001_016+    b_001    tia_h_in_001_016+    1198058.551420872
Rb_h001_016-    b_001    tia_h_in_001_016-    162999.21463987022
Rb_h001_017+    b_001    tia_h_in_001_017+    1198080.8866649424
Rb_h001_017-    b_001    tia_h_in_001_017-    253019.09795351798
Rb_h001_018+    b_001    tia_h_in_001_018+    125615.55560061676
Rb_h001_018-    b_001    tia_h_in_001_018-    1196154.4224094704
Rb_h001_019+    b_001    tia_h_in_001_019+    1196962.9429024728
Rb_h001_019-    b_001    tia_h_in_001_019-    68174.71799375571
Rb_h001_020+    b_001    tia_h_in_001_020+    128664.01337150535
Rb_h001_020-    b_001    tia_h_in_001_020-    1200493.474597998

* ----- Weights
* Layer 002

* Neuron 1
Rh002_001_001+    hidden_activ_out_h001_001    tia_h_in_002_001+    1217409.730551798
Rh002_001_001-    hidden_activ_out_h001_001    tia_h_in_002_001-    29441.557412937975
Rh002_002_001+    hidden_activ_out_h001_002    tia_h_in_002_001+    111108.59240058673
Rh002_002_001-    hidden_activ_out_h001_002    tia_h_in_002_001-    1198135.0993435082
Rh002_003_001+    hidden_activ_out_h001_003    tia_h_in_002_001+    1193439.5662438767
Rh002_003_001-    hidden_activ_out_h001_003    tia_h_in_002_001-    30084.156623847743
Rh002_004_001+    hidden_activ_out_h001_004    tia_h_in_002_001+    1209282.1215619189
Rh002_004_001-    hidden_activ_out_h001_004    tia_h_in_002_001-    1082898.8407583535
Rh002_005_001+    hidden_activ_out_h001_005    tia_h_in_002_001+    20300.42947066616
Rh002_005_001-    hidden_activ_out_h001_005    tia_h_in_002_001-    1193889.9692180476
Rh002_006_001+    hidden_activ_out_h001_006    tia_h_in_002_001+    226267.61725520884
Rh002_006_001-    hidden_activ_out_h001_006    tia_h_in_002_001-    1198824.6782702145
Rh002_007_001+    hidden_activ_out_h001_007    tia_h_in_002_001+    76988.2121133473
Rh002_007_001-    hidden_activ_out_h001_007    tia_h_in_002_001-    1191633.1863401968
Rh002_008_001+    hidden_activ_out_h001_008    tia_h_in_002_001+    21560.89668755685
Rh002_008_001-    hidden_activ_out_h001_008    tia_h_in_002_001-    1208073.2136920267
Rh002_009_001+    hidden_activ_out_h001_009    tia_h_in_002_001+    60568.001332543674
Rh002_009_001-    hidden_activ_out_h001_009    tia_h_in_002_001-    1192836.4672487304
Rh002_010_001+    hidden_activ_out_h001_010    tia_h_in_002_001+    295531.64115768764
Rh002_010_001-    hidden_activ_out_h001_010    tia_h_in_002_001-    1190406.0333051374
Rh002_011_001+    hidden_activ_out_h001_011    tia_h_in_002_001+    38047.21005808193
Rh002_011_001-    hidden_activ_out_h001_011    tia_h_in_002_001-    1189588.282367658
Rh002_012_001+    hidden_activ_out_h001_012    tia_h_in_002_001+    932079.2426228051
Rh002_012_001-    hidden_activ_out_h001_012    tia_h_in_002_001-    1203239.0498891824
Rh002_013_001+    hidden_activ_out_h001_013    tia_h_in_002_001+    38391.683152395075
Rh002_013_001-    hidden_activ_out_h001_013    tia_h_in_002_001-    1200642.594146995
Rh002_014_001+    hidden_activ_out_h001_014    tia_h_in_002_001+    220759.24393744202
Rh002_014_001-    hidden_activ_out_h001_014    tia_h_in_002_001-    1198403.4286912058
Rh002_015_001+    hidden_activ_out_h001_015    tia_h_in_002_001+    1204015.1661989668
Rh002_015_001-    hidden_activ_out_h001_015    tia_h_in_002_001-    798395.5276366443
Rh002_016_001+    hidden_activ_out_h001_016    tia_h_in_002_001+    1204621.0160297912
Rh002_016_001-    hidden_activ_out_h001_016    tia_h_in_002_001-    36010.54335822509
Rh002_017_001+    hidden_activ_out_h001_017    tia_h_in_002_001+    1200399.4469593866
Rh002_017_001-    hidden_activ_out_h001_017    tia_h_in_002_001-    31112.66930068005
Rh002_018_001+    hidden_activ_out_h001_018    tia_h_in_002_001+    85043.11921345771
Rh002_018_001-    hidden_activ_out_h001_018    tia_h_in_002_001-    1227348.1890819531
Rh002_019_001+    hidden_activ_out_h001_019    tia_h_in_002_001+    1214849.6527715183
Rh002_019_001-    hidden_activ_out_h001_019    tia_h_in_002_001-    26901.91664483399
Rh002_020_001+    hidden_activ_out_h001_020    tia_h_in_002_001+    1199322.533406946
Rh002_020_001-    hidden_activ_out_h001_020    tia_h_in_002_001-    664771.2355615816

* Neuron 2
Rh002_001_002+    hidden_activ_out_h001_001    tia_h_in_002_002+    1212623.9008805936
Rh002_001_002-    hidden_activ_out_h001_001    tia_h_in_002_002-    221026.15346198474
Rh002_002_002+    hidden_activ_out_h001_002    tia_h_in_002_002+    1212182.72843338
Rh002_002_002-    hidden_activ_out_h001_002    tia_h_in_002_002-    27073.471153849205
Rh002_003_002+    hidden_activ_out_h001_003    tia_h_in_002_002+    55670.85702201937
Rh002_003_002-    hidden_activ_out_h001_003    tia_h_in_002_002-    1195726.261385706
Rh002_004_002+    hidden_activ_out_h001_004    tia_h_in_002_002+    109752.64581842304
Rh002_004_002-    hidden_activ_out_h001_004    tia_h_in_002_002-    1199229.5924281047
Rh002_005_002+    hidden_activ_out_h001_005    tia_h_in_002_002+    1185522.109130853
Rh002_005_002-    hidden_activ_out_h001_005    tia_h_in_002_002-    46230.90851047596
Rh002_006_002+    hidden_activ_out_h001_006    tia_h_in_002_002+    152112.15971103593
Rh002_006_002-    hidden_activ_out_h001_006    tia_h_in_002_002-    1187586.6019537994
Rh002_007_002+    hidden_activ_out_h001_007    tia_h_in_002_002+    1217807.8932540745
Rh002_007_002-    hidden_activ_out_h001_007    tia_h_in_002_002-    39049.11947703369
Rh002_008_002+    hidden_activ_out_h001_008    tia_h_in_002_002+    1209664.1074688674
Rh002_008_002-    hidden_activ_out_h001_008    tia_h_in_002_002-    39761.15836642706
Rh002_009_002+    hidden_activ_out_h001_009    tia_h_in_002_002+    1200319.2530327113
Rh002_009_002-    hidden_activ_out_h001_009    tia_h_in_002_002-    39079.249815266376
Rh002_010_002+    hidden_activ_out_h001_010    tia_h_in_002_002+    117893.81998837148
Rh002_010_002-    hidden_activ_out_h001_010    tia_h_in_002_002-    1208402.6554206773
Rh002_011_002+    hidden_activ_out_h001_011    tia_h_in_002_002+    1208002.158235823
Rh002_011_002-    hidden_activ_out_h001_011    tia_h_in_002_002-    37014.534563435096
Rh002_012_002+    hidden_activ_out_h001_012    tia_h_in_002_002+    1199888.1409459573
Rh002_012_002-    hidden_activ_out_h001_012    tia_h_in_002_002-    86392.65394698872
Rh002_013_002+    hidden_activ_out_h001_013    tia_h_in_002_002+    1196742.7706691208
Rh002_013_002-    hidden_activ_out_h001_013    tia_h_in_002_002-    33594.82297344162
Rh002_014_002+    hidden_activ_out_h001_014    tia_h_in_002_002+    287634.5282489495
Rh002_014_002-    hidden_activ_out_h001_014    tia_h_in_002_002-    1204318.6828909854
Rh002_015_002+    hidden_activ_out_h001_015    tia_h_in_002_002+    102277.79081574215
Rh002_015_002-    hidden_activ_out_h001_015    tia_h_in_002_002-    1187447.970611377
Rh002_016_002+    hidden_activ_out_h001_016    tia_h_in_002_002+    1214727.3928744209
Rh002_016_002-    hidden_activ_out_h001_016    tia_h_in_002_002-    130695.23534680836
Rh002_017_002+    hidden_activ_out_h001_017    tia_h_in_002_002+    189019.31089963007
Rh002_017_002-    hidden_activ_out_h001_017    tia_h_in_002_002-    1201866.511938218
Rh002_018_002+    hidden_activ_out_h001_018    tia_h_in_002_002+    1209885.328216194
Rh002_018_002-    hidden_activ_out_h001_018    tia_h_in_002_002-    31883.697424545004
Rh002_019_002+    hidden_activ_out_h001_019    tia_h_in_002_002+    51548.254948448644
Rh002_019_002-    hidden_activ_out_h001_019    tia_h_in_002_002-    1208152.323470537
Rh002_020_002+    hidden_activ_out_h001_020    tia_h_in_002_002+    1194440.7297127086
Rh002_020_002-    hidden_activ_out_h001_020    tia_h_in_002_002-    46377.2059302316

* Neuron 3
Rh002_001_003+    hidden_activ_out_h001_001    tia_h_in_002_003+    58025.941142189644
Rh002_001_003-    hidden_activ_out_h001_001    tia_h_in_002_003-    1213426.0641412714
Rh002_002_003+    hidden_activ_out_h001_002    tia_h_in_002_003+    1217514.982225307
Rh002_002_003-    hidden_activ_out_h001_002    tia_h_in_002_003-    30150.741703842774
Rh002_003_003+    hidden_activ_out_h001_003    tia_h_in_002_003+    94754.25644941286
Rh002_003_003-    hidden_activ_out_h001_003    tia_h_in_002_003-    1202405.5745875223
Rh002_004_003+    hidden_activ_out_h001_004    tia_h_in_002_003+    159183.10358898563
Rh002_004_003-    hidden_activ_out_h001_004    tia_h_in_002_003-    1188215.226641444
Rh002_005_003+    hidden_activ_out_h001_005    tia_h_in_002_003+    1202854.3770857083
Rh002_005_003-    hidden_activ_out_h001_005    tia_h_in_002_003-    64557.10572983896
Rh002_006_003+    hidden_activ_out_h001_006    tia_h_in_002_003+    275507.7990074949
Rh002_006_003-    hidden_activ_out_h001_006    tia_h_in_002_003-    1197883.9222620348
Rh002_007_003+    hidden_activ_out_h001_007    tia_h_in_002_003+    1203582.1600979
Rh002_007_003-    hidden_activ_out_h001_007    tia_h_in_002_003-    83469.81301297752
Rh002_008_003+    hidden_activ_out_h001_008    tia_h_in_002_003+    1197417.6611777137
Rh002_008_003-    hidden_activ_out_h001_008    tia_h_in_002_003-    105800.02950569653
Rh002_009_003+    hidden_activ_out_h001_009    tia_h_in_002_003+    1203250.004009937
Rh002_009_003-    hidden_activ_out_h001_009    tia_h_in_002_003-    47038.518539890014
Rh002_010_003+    hidden_activ_out_h001_010    tia_h_in_002_003+    205432.14875248377
Rh002_010_003-    hidden_activ_out_h001_010    tia_h_in_002_003-    1208867.0093034352
Rh002_011_003+    hidden_activ_out_h001_011    tia_h_in_002_003+    1204129.6951170252
Rh002_011_003-    hidden_activ_out_h001_011    tia_h_in_002_003-    51395.65244356995
Rh002_012_003+    hidden_activ_out_h001_012    tia_h_in_002_003+    1208849.3747874892
Rh002_012_003-    hidden_activ_out_h001_012    tia_h_in_002_003-    128033.51730241203
Rh002_013_003+    hidden_activ_out_h001_013    tia_h_in_002_003+    1208235.6736860857
Rh002_013_003-    hidden_activ_out_h001_013    tia_h_in_002_003-    45889.99842667496
Rh002_014_003+    hidden_activ_out_h001_014    tia_h_in_002_003+    124492.98787578174
Rh002_014_003-    hidden_activ_out_h001_014    tia_h_in_002_003-    1187042.2001290526
Rh002_015_003+    hidden_activ_out_h001_015    tia_h_in_002_003+    192166.66260310548
Rh002_015_003-    hidden_activ_out_h001_015    tia_h_in_002_003-    1181386.8361883918
Rh002_016_003+    hidden_activ_out_h001_016    tia_h_in_002_003+    61588.842155712
Rh002_016_003-    hidden_activ_out_h001_016    tia_h_in_002_003-    1205598.7641999568
Rh002_017_003+    hidden_activ_out_h001_017    tia_h_in_002_003+    1211691.9371909916
Rh002_017_003-    hidden_activ_out_h001_017    tia_h_in_002_003-    97588.9077754935
Rh002_018_003+    hidden_activ_out_h001_018    tia_h_in_002_003+    1215542.5279198557
Rh002_018_003-    hidden_activ_out_h001_018    tia_h_in_002_003-    92740.97128745902
Rh002_019_003+    hidden_activ_out_h001_019    tia_h_in_002_003+    113931.45930277603
Rh002_019_003-    hidden_activ_out_h001_019    tia_h_in_002_003-    1202881.9337432585
Rh002_020_003+    hidden_activ_out_h001_020    tia_h_in_002_003+    1199011.5330498936
Rh002_020_003-    hidden_activ_out_h001_020    tia_h_in_002_003-    310569.0164893475

* Neuron 4
Rh002_001_004+    hidden_activ_out_h001_001    tia_h_in_002_004+    38971.90947303225
Rh002_001_004-    hidden_activ_out_h001_001    tia_h_in_002_004-    1194203.6015893437
Rh002_002_004+    hidden_activ_out_h001_002    tia_h_in_002_004+    1212058.2686338928
Rh002_002_004-    hidden_activ_out_h001_002    tia_h_in_002_004-    119756.7182723278
Rh002_003_004+    hidden_activ_out_h001_003    tia_h_in_002_004+    68432.21026835087
Rh002_003_004-    hidden_activ_out_h001_003    tia_h_in_002_004-    1188161.2028585188
Rh002_004_004+    hidden_activ_out_h001_004    tia_h_in_002_004+    1204427.6576516968
Rh002_004_004-    hidden_activ_out_h001_004    tia_h_in_002_004-    930306.1992039469
Rh002_005_004+    hidden_activ_out_h001_005    tia_h_in_002_004+    1188903.278612401
Rh002_005_004-    hidden_activ_out_h001_005    tia_h_in_002_004-    83536.55906843035
Rh002_006_004+    hidden_activ_out_h001_006    tia_h_in_002_004+    110646.39213000759
Rh002_006_004-    hidden_activ_out_h001_006    tia_h_in_002_004-    1197755.0714585932
Rh002_007_004+    hidden_activ_out_h001_007    tia_h_in_002_004+    1208619.8543885658
Rh002_007_004-    hidden_activ_out_h001_007    tia_h_in_002_004-    181567.05121638012
Rh002_008_004+    hidden_activ_out_h001_008    tia_h_in_002_004+    1206581.2253120446
Rh002_008_004-    hidden_activ_out_h001_008    tia_h_in_002_004-    124649.71713238343
Rh002_009_004+    hidden_activ_out_h001_009    tia_h_in_002_004+    436287.4646155273
Rh002_009_004-    hidden_activ_out_h001_009    tia_h_in_002_004-    1197720.866277313
Rh002_010_004+    hidden_activ_out_h001_010    tia_h_in_002_004+    1195350.126253259
Rh002_010_004-    hidden_activ_out_h001_010    tia_h_in_002_004-    479862.6028011797
Rh002_011_004+    hidden_activ_out_h001_011    tia_h_in_002_004+    1205099.7136019159
Rh002_011_004-    hidden_activ_out_h001_011    tia_h_in_002_004-    187241.15509031605
Rh002_012_004+    hidden_activ_out_h001_012    tia_h_in_002_004+    410931.0070457669
Rh002_012_004-    hidden_activ_out_h001_012    tia_h_in_002_004-    1211143.6774373017
Rh002_013_004+    hidden_activ_out_h001_013    tia_h_in_002_004+    1194510.4199662602
Rh002_013_004-    hidden_activ_out_h001_013    tia_h_in_002_004-    276782.2848133737
Rh002_014_004+    hidden_activ_out_h001_014    tia_h_in_002_004+    317074.8821960531
Rh002_014_004-    hidden_activ_out_h001_014    tia_h_in_002_004-    1195022.340666443
Rh002_015_004+    hidden_activ_out_h001_015    tia_h_in_002_004+    117834.93628571306
Rh002_015_004-    hidden_activ_out_h001_015    tia_h_in_002_004-    1186181.8508346865
Rh002_016_004+    hidden_activ_out_h001_016    tia_h_in_002_004+    41398.64105250329
Rh002_016_004-    hidden_activ_out_h001_016    tia_h_in_002_004-    1200675.499573237
Rh002_017_004+    hidden_activ_out_h001_017    tia_h_in_002_004+    58873.517827144555
Rh002_017_004-    hidden_activ_out_h001_017    tia_h_in_002_004-    1193209.5232024638
Rh002_018_004+    hidden_activ_out_h001_018    tia_h_in_002_004+    351962.8999001081
Rh002_018_004-    hidden_activ_out_h001_018    tia_h_in_002_004-    1183823.7054071533
Rh002_019_004+    hidden_activ_out_h001_019    tia_h_in_002_004+    48194.95856809881
Rh002_019_004-    hidden_activ_out_h001_019    tia_h_in_002_004-    1205718.475251194
Rh002_020_004+    hidden_activ_out_h001_020    tia_h_in_002_004+    252316.6317008808
Rh002_020_004-    hidden_activ_out_h001_020    tia_h_in_002_004-    1200709.385320639

* Neuron 5
Rh002_001_005+    hidden_activ_out_h001_001    tia_h_in_002_005+    48848.15442011114
Rh002_001_005-    hidden_activ_out_h001_001    tia_h_in_002_005-    1209542.0808965806
Rh002_002_005+    hidden_activ_out_h001_002    tia_h_in_002_005+    1211142.0909223268
Rh002_002_005-    hidden_activ_out_h001_002    tia_h_in_002_005-    108599.02614799888
Rh002_003_005+    hidden_activ_out_h001_003    tia_h_in_002_005+    82596.40735676231
Rh002_003_005-    hidden_activ_out_h001_003    tia_h_in_002_005-    1197609.6810701406
Rh002_004_005+    hidden_activ_out_h001_004    tia_h_in_002_005+    167438.61841008073
Rh002_004_005-    hidden_activ_out_h001_004    tia_h_in_002_005-    1193375.7451032903
Rh002_005_005+    hidden_activ_out_h001_005    tia_h_in_002_005+    1196797.4019327841
Rh002_005_005-    hidden_activ_out_h001_005    tia_h_in_002_005-    63799.29872163788
Rh002_006_005+    hidden_activ_out_h001_006    tia_h_in_002_005+    1197460.077651902
Rh002_006_005-    hidden_activ_out_h001_006    tia_h_in_002_005-    519069.2319742487
Rh002_007_005+    hidden_activ_out_h001_007    tia_h_in_002_005+    1202158.0424593955
Rh002_007_005-    hidden_activ_out_h001_007    tia_h_in_002_005-    174419.2663385638
Rh002_008_005+    hidden_activ_out_h001_008    tia_h_in_002_005+    1197210.5485503355
Rh002_008_005-    hidden_activ_out_h001_008    tia_h_in_002_005-    110920.00892903586
Rh002_009_005+    hidden_activ_out_h001_009    tia_h_in_002_005+    1204358.878809586
Rh002_009_005-    hidden_activ_out_h001_009    tia_h_in_002_005-    870897.1788574985
Rh002_010_005+    hidden_activ_out_h001_010    tia_h_in_002_005+    337035.02231423714
Rh002_010_005-    hidden_activ_out_h001_010    tia_h_in_002_005-    1216047.0577105626
Rh002_011_005+    hidden_activ_out_h001_011    tia_h_in_002_005+    1200918.2419991056
Rh002_011_005-    hidden_activ_out_h001_011    tia_h_in_002_005-    151527.5962603411
Rh002_012_005+    hidden_activ_out_h001_012    tia_h_in_002_005+    312732.9567567917
Rh002_012_005-    hidden_activ_out_h001_012    tia_h_in_002_005-    1198106.7498082933
Rh002_013_005+    hidden_activ_out_h001_013    tia_h_in_002_005+    1191884.5172592278
Rh002_013_005-    hidden_activ_out_h001_013    tia_h_in_002_005-    228153.12353385793
Rh002_014_005+    hidden_activ_out_h001_014    tia_h_in_002_005+    188678.02090747916
Rh002_014_005-    hidden_activ_out_h001_014    tia_h_in_002_005-    1211971.1478811305
Rh002_015_005+    hidden_activ_out_h001_015    tia_h_in_002_005+    1049169.0586420828
Rh002_015_005-    hidden_activ_out_h001_015    tia_h_in_002_005-    1220966.7614337844
Rh002_016_005+    hidden_activ_out_h001_016    tia_h_in_002_005+    51310.767680983015
Rh002_016_005-    hidden_activ_out_h001_016    tia_h_in_002_005-    1205595.8152027773
Rh002_017_005+    hidden_activ_out_h001_017    tia_h_in_002_005+    77940.65648337411
Rh002_017_005-    hidden_activ_out_h001_017    tia_h_in_002_005-    1180006.7818101353
Rh002_018_005+    hidden_activ_out_h001_018    tia_h_in_002_005+    374476.9870599533
Rh002_018_005-    hidden_activ_out_h001_018    tia_h_in_002_005-    1203808.5119064073
Rh002_019_005+    hidden_activ_out_h001_019    tia_h_in_002_005+    60463.90284353736
Rh002_019_005-    hidden_activ_out_h001_019    tia_h_in_002_005-    1195125.3070546575
Rh002_020_005+    hidden_activ_out_h001_020    tia_h_in_002_005+    187616.08975100107
Rh002_020_005-    hidden_activ_out_h001_020    tia_h_in_002_005-    1194880.3038884022

* Neuron 6
Rh002_001_006+    hidden_activ_out_h001_001    tia_h_in_002_006+    1191163.8244648818
Rh002_001_006-    hidden_activ_out_h001_001    tia_h_in_002_006-    26884.70598044434
Rh002_002_006+    hidden_activ_out_h001_002    tia_h_in_002_006+    111634.74162588354
Rh002_002_006-    hidden_activ_out_h001_002    tia_h_in_002_006-    1192900.3843858514
Rh002_003_006+    hidden_activ_out_h001_003    tia_h_in_002_006+    1218228.8276864558
Rh002_003_006-    hidden_activ_out_h001_003    tia_h_in_002_006-    23588.898060503852
Rh002_004_006+    hidden_activ_out_h001_004    tia_h_in_002_006+    237918.1404354604
Rh002_004_006-    hidden_activ_out_h001_004    tia_h_in_002_006-    1193145.8258948796
Rh002_005_006+    hidden_activ_out_h001_005    tia_h_in_002_006+    22427.797445042364
Rh002_005_006-    hidden_activ_out_h001_005    tia_h_in_002_006-    1192581.6583817967
Rh002_006_006+    hidden_activ_out_h001_006    tia_h_in_002_006+    197541.3750961745
Rh002_006_006-    hidden_activ_out_h001_006    tia_h_in_002_006-    1201761.6126721702
Rh002_007_006+    hidden_activ_out_h001_007    tia_h_in_002_006+    74227.77760420243
Rh002_007_006-    hidden_activ_out_h001_007    tia_h_in_002_006-    1198470.4547679618
Rh002_008_006+    hidden_activ_out_h001_008    tia_h_in_002_006+    26408.8935646162
Rh002_008_006-    hidden_activ_out_h001_008    tia_h_in_002_006-    1194210.6746004717
Rh002_009_006+    hidden_activ_out_h001_009    tia_h_in_002_006+    82570.56558582374
Rh002_009_006-    hidden_activ_out_h001_009    tia_h_in_002_006-    1202883.3757981672
Rh002_010_006+    hidden_activ_out_h001_010    tia_h_in_002_006+    542275.3040137134
Rh002_010_006-    hidden_activ_out_h001_010    tia_h_in_002_006-    1205880.7087831784
Rh002_011_006+    hidden_activ_out_h001_011    tia_h_in_002_006+    47304.618998487735
Rh002_011_006-    hidden_activ_out_h001_011    tia_h_in_002_006-    1203501.6846783678
Rh002_012_006+    hidden_activ_out_h001_012    tia_h_in_002_006+    399454.96766624064
Rh002_012_006-    hidden_activ_out_h001_012    tia_h_in_002_006-    1188881.458926506
Rh002_013_006+    hidden_activ_out_h001_013    tia_h_in_002_006+    46361.504650238116
Rh002_013_006-    hidden_activ_out_h001_013    tia_h_in_002_006-    1202571.7095610206
Rh002_014_006+    hidden_activ_out_h001_014    tia_h_in_002_006+    179821.52968546972
Rh002_014_006-    hidden_activ_out_h001_014    tia_h_in_002_006-    1193648.4556011115
Rh002_015_006+    hidden_activ_out_h001_015    tia_h_in_002_006+    226841.42034380822
Rh002_015_006-    hidden_activ_out_h001_015    tia_h_in_002_006-    1192451.119447387
Rh002_016_006+    hidden_activ_out_h001_016    tia_h_in_002_006+    1178687.7292785957
Rh002_016_006-    hidden_activ_out_h001_016    tia_h_in_002_006-    31200.822921240324
Rh002_017_006+    hidden_activ_out_h001_017    tia_h_in_002_006+    1210010.23991018
Rh002_017_006-    hidden_activ_out_h001_017    tia_h_in_002_006-    57821.808963553936
Rh002_018_006+    hidden_activ_out_h001_018    tia_h_in_002_006+    58099.93331975444
Rh002_018_006-    hidden_activ_out_h001_018    tia_h_in_002_006-    1204325.922626812
Rh002_019_006+    hidden_activ_out_h001_019    tia_h_in_002_006+    1199933.871656285
Rh002_019_006-    hidden_activ_out_h001_019    tia_h_in_002_006-    20071.816866650002
Rh002_020_006+    hidden_activ_out_h001_020    tia_h_in_002_006+    1207321.9161364771
Rh002_020_006-    hidden_activ_out_h001_020    tia_h_in_002_006-    521979.5987501605

* Neuron 7
Rh002_001_007+    hidden_activ_out_h001_001    tia_h_in_002_007+    80556.4706521557
Rh002_001_007-    hidden_activ_out_h001_001    tia_h_in_002_007-    1189646.1135580211
Rh002_002_007+    hidden_activ_out_h001_002    tia_h_in_002_007+    1193519.6802688497
Rh002_002_007-    hidden_activ_out_h001_002    tia_h_in_002_007-    40551.87796244787
Rh002_003_007+    hidden_activ_out_h001_003    tia_h_in_002_007+    63262.4613788448
Rh002_003_007-    hidden_activ_out_h001_003    tia_h_in_002_007-    1207634.0845002201
Rh002_004_007+    hidden_activ_out_h001_004    tia_h_in_002_007+    347493.19944297237
Rh002_004_007-    hidden_activ_out_h001_004    tia_h_in_002_007-    1200950.545413693
Rh002_005_007+    hidden_activ_out_h001_005    tia_h_in_002_007+    1200103.8012384768
Rh002_005_007-    hidden_activ_out_h001_005    tia_h_in_002_007-    44002.633778826435
Rh002_006_007+    hidden_activ_out_h001_006    tia_h_in_002_007+    381058.9599134128
Rh002_006_007-    hidden_activ_out_h001_006    tia_h_in_002_007-    1189280.9472430982
Rh002_007_007+    hidden_activ_out_h001_007    tia_h_in_002_007+    1196160.3971252488
Rh002_007_007-    hidden_activ_out_h001_007    tia_h_in_002_007-    73320.25590580562
Rh002_008_007+    hidden_activ_out_h001_008    tia_h_in_002_007+    1192786.9173164351
Rh002_008_007-    hidden_activ_out_h001_008    tia_h_in_002_007-    100312.91581549088
Rh002_009_007+    hidden_activ_out_h001_009    tia_h_in_002_007+    1183034.0318501294
Rh002_009_007-    hidden_activ_out_h001_009    tia_h_in_002_007-    73943.71715148867
Rh002_010_007+    hidden_activ_out_h001_010    tia_h_in_002_007+    104060.9120973098
Rh002_010_007-    hidden_activ_out_h001_010    tia_h_in_002_007-    1193579.6797513047
Rh002_011_007+    hidden_activ_out_h001_011    tia_h_in_002_007+    1203423.1815112715
Rh002_011_007-    hidden_activ_out_h001_011    tia_h_in_002_007-    56197.05254528644
Rh002_012_007+    hidden_activ_out_h001_012    tia_h_in_002_007+    1203450.9050967775
Rh002_012_007-    hidden_activ_out_h001_012    tia_h_in_002_007-    235912.8922949481
Rh002_013_007+    hidden_activ_out_h001_013    tia_h_in_002_007+    1189754.3259092937
Rh002_013_007-    hidden_activ_out_h001_013    tia_h_in_002_007-    48984.79900106932
Rh002_014_007+    hidden_activ_out_h001_014    tia_h_in_002_007+    127990.22212195267
Rh002_014_007-    hidden_activ_out_h001_014    tia_h_in_002_007-    1200592.7700930722
Rh002_015_007+    hidden_activ_out_h001_015    tia_h_in_002_007+    1204377.4320955705
Rh002_015_007-    hidden_activ_out_h001_015    tia_h_in_002_007-    773429.0415604259
Rh002_016_007+    hidden_activ_out_h001_016    tia_h_in_002_007+    67609.91727749007
Rh002_016_007-    hidden_activ_out_h001_016    tia_h_in_002_007-    1212679.2175518256
Rh002_017_007+    hidden_activ_out_h001_017    tia_h_in_002_007+    179652.9654084976
Rh002_017_007-    hidden_activ_out_h001_017    tia_h_in_002_007-    1197879.2867049929
Rh002_018_007+    hidden_activ_out_h001_018    tia_h_in_002_007+    1183113.280671651
Rh002_018_007-    hidden_activ_out_h001_018    tia_h_in_002_007-    164280.2277635492
Rh002_019_007+    hidden_activ_out_h001_019    tia_h_in_002_007+    63228.786190589686
Rh002_019_007-    hidden_activ_out_h001_019    tia_h_in_002_007-    1198861.2055644111
Rh002_020_007+    hidden_activ_out_h001_020    tia_h_in_002_007+    680660.5373029173
Rh002_020_007-    hidden_activ_out_h001_020    tia_h_in_002_007-    1198353.6770526238

* Neuron 8
Rh002_001_008+    hidden_activ_out_h001_001    tia_h_in_002_008+    186157.7212208313
Rh002_001_008-    hidden_activ_out_h001_001    tia_h_in_002_008-    1194573.6392448551
Rh002_002_008+    hidden_activ_out_h001_002    tia_h_in_002_008+    1202211.0890967303
Rh002_002_008-    hidden_activ_out_h001_002    tia_h_in_002_008-    22143.958985618592
Rh002_003_008+    hidden_activ_out_h001_003    tia_h_in_002_008+    71552.1091974911
Rh002_003_008-    hidden_activ_out_h001_003    tia_h_in_002_008-    1188248.1058100064
Rh002_004_008+    hidden_activ_out_h001_004    tia_h_in_002_008+    147419.11160960852
Rh002_004_008-    hidden_activ_out_h001_004    tia_h_in_002_008-    1199324.8092302938
Rh002_005_008+    hidden_activ_out_h001_005    tia_h_in_002_008+    1186763.4621503172
Rh002_005_008-    hidden_activ_out_h001_005    tia_h_in_002_008-    53137.282764994925
Rh002_006_008+    hidden_activ_out_h001_006    tia_h_in_002_008+    418612.3488653932
Rh002_006_008-    hidden_activ_out_h001_006    tia_h_in_002_008-    1197403.827716035
Rh002_007_008+    hidden_activ_out_h001_007    tia_h_in_002_008+    1192143.790225106
Rh002_007_008-    hidden_activ_out_h001_007    tia_h_in_002_008-    39099.899437310116
Rh002_008_008+    hidden_activ_out_h001_008    tia_h_in_002_008+    1185436.1051270608
Rh002_008_008-    hidden_activ_out_h001_008    tia_h_in_002_008-    55457.83484472165
Rh002_009_008+    hidden_activ_out_h001_009    tia_h_in_002_008+    1206872.7864522114
Rh002_009_008-    hidden_activ_out_h001_009    tia_h_in_002_008-    28732.621486812837
Rh002_010_008+    hidden_activ_out_h001_010    tia_h_in_002_008+    104713.7811726721
Rh002_010_008-    hidden_activ_out_h001_010    tia_h_in_002_008-    1193559.0182398448
Rh002_011_008+    hidden_activ_out_h001_011    tia_h_in_002_008+    1199483.497588185
Rh002_011_008-    hidden_activ_out_h001_011    tia_h_in_002_008-    51217.777261716095
Rh002_012_008+    hidden_activ_out_h001_012    tia_h_in_002_008+    1208963.1989445314
Rh002_012_008-    hidden_activ_out_h001_012    tia_h_in_002_008-    51904.249191874835
Rh002_013_008+    hidden_activ_out_h001_013    tia_h_in_002_008+    1211872.338597773
Rh002_013_008-    hidden_activ_out_h001_013    tia_h_in_002_008-    35288.212776846354
Rh002_014_008+    hidden_activ_out_h001_014    tia_h_in_002_008+    163753.24687682965
Rh002_014_008-    hidden_activ_out_h001_014    tia_h_in_002_008-    1190291.9346461322
Rh002_015_008+    hidden_activ_out_h001_015    tia_h_in_002_008+    116446.27281762747
Rh002_015_008-    hidden_activ_out_h001_015    tia_h_in_002_008-    1198822.8866252191
Rh002_016_008+    hidden_activ_out_h001_016    tia_h_in_002_008+    243285.23076503235
Rh002_016_008-    hidden_activ_out_h001_016    tia_h_in_002_008-    1191732.8910870105
Rh002_017_008+    hidden_activ_out_h001_017    tia_h_in_002_008+    1189911.0565528336
Rh002_017_008-    hidden_activ_out_h001_017    tia_h_in_002_008-    265909.68264204916
Rh002_018_008+    hidden_activ_out_h001_018    tia_h_in_002_008+    1199083.2943745146
Rh002_018_008-    hidden_activ_out_h001_018    tia_h_in_002_008-    26378.11564824194
Rh002_019_008+    hidden_activ_out_h001_019    tia_h_in_002_008+    75704.70156563689
Rh002_019_008-    hidden_activ_out_h001_019    tia_h_in_002_008-    1191845.9474262586
Rh002_020_008+    hidden_activ_out_h001_020    tia_h_in_002_008+    1217486.5347523957
Rh002_020_008-    hidden_activ_out_h001_020    tia_h_in_002_008-    29328.50125481534

* Neuron 9
Rh002_001_009+    hidden_activ_out_h001_001    tia_h_in_002_009+    207665.10062064114
Rh002_001_009-    hidden_activ_out_h001_001    tia_h_in_002_009-    1200929.2935482888
Rh002_002_009+    hidden_activ_out_h001_002    tia_h_in_002_009+    1204776.242847943
Rh002_002_009-    hidden_activ_out_h001_002    tia_h_in_002_009-    35038.885062132904
Rh002_003_009+    hidden_activ_out_h001_003    tia_h_in_002_009+    53370.90245344495
Rh002_003_009-    hidden_activ_out_h001_003    tia_h_in_002_009-    1187630.1190286037
Rh002_004_009+    hidden_activ_out_h001_004    tia_h_in_002_009+    285524.45728458016
Rh002_004_009-    hidden_activ_out_h001_004    tia_h_in_002_009-    1196681.5306782897
Rh002_005_009+    hidden_activ_out_h001_005    tia_h_in_002_009+    1192615.6473070362
Rh002_005_009-    hidden_activ_out_h001_005    tia_h_in_002_009-    42391.89328900563
Rh002_006_009+    hidden_activ_out_h001_006    tia_h_in_002_009+    108781.98933554832
Rh002_006_009-    hidden_activ_out_h001_006    tia_h_in_002_009-    1198366.7598187842
Rh002_007_009+    hidden_activ_out_h001_007    tia_h_in_002_009+    1202758.1666134186
Rh002_007_009-    hidden_activ_out_h001_007    tia_h_in_002_009-    53977.831301559854
Rh002_008_009+    hidden_activ_out_h001_008    tia_h_in_002_009+    1200057.7361316083
Rh002_008_009-    hidden_activ_out_h001_008    tia_h_in_002_009-    57068.40568533497
Rh002_009_009+    hidden_activ_out_h001_009    tia_h_in_002_009+    1209837.100177836
Rh002_009_009-    hidden_activ_out_h001_009    tia_h_in_002_009-    36789.02087168468
Rh002_010_009+    hidden_activ_out_h001_010    tia_h_in_002_009+    121137.28315754519
Rh002_010_009-    hidden_activ_out_h001_010    tia_h_in_002_009-    1205276.318511714
Rh002_011_009+    hidden_activ_out_h001_011    tia_h_in_002_009+    1208478.5650030435
Rh002_011_009-    hidden_activ_out_h001_011    tia_h_in_002_009-    46454.77981210603
Rh002_012_009+    hidden_activ_out_h001_012    tia_h_in_002_009+    1193298.2322312666
Rh002_012_009-    hidden_activ_out_h001_012    tia_h_in_002_009-    103733.01661746878
Rh002_013_009+    hidden_activ_out_h001_013    tia_h_in_002_009+    1200298.810499077
Rh002_013_009-    hidden_activ_out_h001_013    tia_h_in_002_009-    32407.158926446435
Rh002_014_009+    hidden_activ_out_h001_014    tia_h_in_002_009+    150294.4537804259
Rh002_014_009-    hidden_activ_out_h001_014    tia_h_in_002_009-    1205399.2583348006
Rh002_015_009+    hidden_activ_out_h001_015    tia_h_in_002_009+    227839.2218346612
Rh002_015_009-    hidden_activ_out_h001_015    tia_h_in_002_009-    1201775.0859436847
Rh002_016_009+    hidden_activ_out_h001_016    tia_h_in_002_009+    276558.715480429
Rh002_016_009-    hidden_activ_out_h001_016    tia_h_in_002_009-    1191932.7244577685
Rh002_017_009+    hidden_activ_out_h001_017    tia_h_in_002_009+    255386.88373183928
Rh002_017_009-    hidden_activ_out_h001_017    tia_h_in_002_009-    1183284.0381158742
Rh002_018_009+    hidden_activ_out_h001_018    tia_h_in_002_009+    1193074.5262350636
Rh002_018_009-    hidden_activ_out_h001_018    tia_h_in_002_009-    61527.28068961589
Rh002_019_009+    hidden_activ_out_h001_019    tia_h_in_002_009+    72943.33647723144
Rh002_019_009-    hidden_activ_out_h001_019    tia_h_in_002_009-    1210771.5306094852
Rh002_020_009+    hidden_activ_out_h001_020    tia_h_in_002_009+    1202402.4618123882
Rh002_020_009-    hidden_activ_out_h001_020    tia_h_in_002_009-    229664.88319343486

* Neuron 10
Rh002_001_010+    hidden_activ_out_h001_001    tia_h_in_002_010+    44835.178625760076
Rh002_001_010-    hidden_activ_out_h001_001    tia_h_in_002_010-    1196062.617351614
Rh002_002_010+    hidden_activ_out_h001_002    tia_h_in_002_010+    1203773.3112346435
Rh002_002_010-    hidden_activ_out_h001_002    tia_h_in_002_010-    124853.00775566633
Rh002_003_010+    hidden_activ_out_h001_003    tia_h_in_002_010+    59949.130163017435
Rh002_003_010-    hidden_activ_out_h001_003    tia_h_in_002_010-    1202135.7790589123
Rh002_004_010+    hidden_activ_out_h001_004    tia_h_in_002_010+    127800.1833053708
Rh002_004_010-    hidden_activ_out_h001_004    tia_h_in_002_010-    1199343.293162973
Rh002_005_010+    hidden_activ_out_h001_005    tia_h_in_002_010+    1202015.8905596375
Rh002_005_010-    hidden_activ_out_h001_005    tia_h_in_002_010-    71645.2718996233
Rh002_006_010+    hidden_activ_out_h001_006    tia_h_in_002_010+    105162.12519069888
Rh002_006_010-    hidden_activ_out_h001_006    tia_h_in_002_010-    1206210.3682347033
Rh002_007_010+    hidden_activ_out_h001_007    tia_h_in_002_010+    1196972.1536517912
Rh002_007_010-    hidden_activ_out_h001_007    tia_h_in_002_010-    160967.75550499186
Rh002_008_010+    hidden_activ_out_h001_008    tia_h_in_002_010+    1201493.7676563489
Rh002_008_010-    hidden_activ_out_h001_008    tia_h_in_002_010-    93310.76385280519
Rh002_009_010+    hidden_activ_out_h001_009    tia_h_in_002_010+    1192813.0936287562
Rh002_009_010-    hidden_activ_out_h001_009    tia_h_in_002_010-    581635.0010040585
Rh002_010_010+    hidden_activ_out_h001_010    tia_h_in_002_010+    947475.0321700254
Rh002_010_010-    hidden_activ_out_h001_010    tia_h_in_002_010-    1205621.4603178005
Rh002_011_010+    hidden_activ_out_h001_011    tia_h_in_002_010+    1201849.194576022
Rh002_011_010-    hidden_activ_out_h001_011    tia_h_in_002_010-    161108.7190016101
Rh002_012_010+    hidden_activ_out_h001_012    tia_h_in_002_010+    340790.0701420063
Rh002_012_010-    hidden_activ_out_h001_012    tia_h_in_002_010-    1201817.4091874766
Rh002_013_010+    hidden_activ_out_h001_013    tia_h_in_002_010+    1211206.2653414696
Rh002_013_010-    hidden_activ_out_h001_013    tia_h_in_002_010-    249163.57408330878
Rh002_014_010+    hidden_activ_out_h001_014    tia_h_in_002_010+    196550.1285563392
Rh002_014_010-    hidden_activ_out_h001_014    tia_h_in_002_010-    1213660.400419528
Rh002_015_010+    hidden_activ_out_h001_015    tia_h_in_002_010+    132930.14385254707
Rh002_015_010-    hidden_activ_out_h001_015    tia_h_in_002_010-    1209161.4025288085
Rh002_016_010+    hidden_activ_out_h001_016    tia_h_in_002_010+    44157.85162392379
Rh002_016_010-    hidden_activ_out_h001_016    tia_h_in_002_010-    1194203.568775287
Rh002_017_010+    hidden_activ_out_h001_017    tia_h_in_002_010+    67502.65133690648
Rh002_017_010-    hidden_activ_out_h001_017    tia_h_in_002_010-    1204881.0193775396
Rh002_018_010+    hidden_activ_out_h001_018    tia_h_in_002_010+    384299.6781616611
Rh002_018_010-    hidden_activ_out_h001_018    tia_h_in_002_010-    1199716.2367781363
Rh002_019_010+    hidden_activ_out_h001_019    tia_h_in_002_010+    57331.40723972208
Rh002_019_010-    hidden_activ_out_h001_019    tia_h_in_002_010-    1193141.3792660462
Rh002_020_010+    hidden_activ_out_h001_020    tia_h_in_002_010+    202822.45790215337
Rh002_020_010-    hidden_activ_out_h001_020    tia_h_in_002_010-    1208314.3423759784

* ----- Bias
    
        
Rb_h002_001+    b_002    tia_h_in_002_001+    213444.0455082236
Rb_h002_001-    b_002    tia_h_in_002_001-    1199104.5198619524
Rb_h002_002+    b_002    tia_h_in_002_002+    157294.49647853797
Rb_h002_002-    b_002    tia_h_in_002_002-    1179056.0480314633
Rb_h002_003+    b_002    tia_h_in_002_003+    138211.39605232966
Rb_h002_003-    b_002    tia_h_in_002_003-    1213414.5048488735
Rb_h002_004+    b_002    tia_h_in_002_004+    345877.9445413361
Rb_h002_004-    b_002    tia_h_in_002_004-    1198634.3529216505
Rb_h002_005+    b_002    tia_h_in_002_005+    345850.05160424043
Rb_h002_005-    b_002    tia_h_in_002_005-    1211431.6934211354
Rb_h002_006+    b_002    tia_h_in_002_006+    215691.9978823526
Rb_h002_006-    b_002    tia_h_in_002_006-    1191966.6368757316
Rb_h002_007+    b_002    tia_h_in_002_007+    151945.04072365834
Rb_h002_007-    b_002    tia_h_in_002_007-    1207174.2977574193
Rb_h002_008+    b_002    tia_h_in_002_008+    116059.1482238172
Rb_h002_008-    b_002    tia_h_in_002_008-    1206245.6939133396
Rb_h002_009+    b_002    tia_h_in_002_009+    125625.41598474467
Rb_h002_009-    b_002    tia_h_in_002_009-    1197250.2257253474
Rb_h002_010+    b_002    tia_h_in_002_010+    333449.49114257726
Rb_h002_010-    b_002    tia_h_in_002_010-    1216335.8358391207

* ----- Weights
* Layer 003

* Neuron 1
Rh003_001_001+    hidden_activ_out_h002_001    tia_h_in_003_001+    1198293.4118674635
Rh003_001_001-    hidden_activ_out_h002_001    tia_h_in_003_001-    20623.837694179718
Rh003_002_001+    hidden_activ_out_h002_002    tia_h_in_003_001+    20310.520769511637
Rh003_002_001-    hidden_activ_out_h002_002    tia_h_in_003_001-    1198620.8042020178
Rh003_003_001+    hidden_activ_out_h002_003    tia_h_in_003_001+    32305.377684172425
Rh003_003_001-    hidden_activ_out_h002_003    tia_h_in_003_001-    1184979.215835261
Rh003_004_001+    hidden_activ_out_h002_004    tia_h_in_003_001+    69241.9065391741
Rh003_004_001-    hidden_activ_out_h002_004    tia_h_in_003_001-    1217230.0225714846
Rh003_005_001+    hidden_activ_out_h002_005    tia_h_in_003_001+    50839.81234470057
Rh003_005_001-    hidden_activ_out_h002_005    tia_h_in_003_001-    1198881.5549319992
Rh003_006_001+    hidden_activ_out_h002_006    tia_h_in_003_001+    1196017.8220470536
Rh003_006_001-    hidden_activ_out_h002_006    tia_h_in_003_001-    20230.56910790058
Rh003_007_001+    hidden_activ_out_h002_007    tia_h_in_003_001+    40105.580102769985
Rh003_007_001-    hidden_activ_out_h002_007    tia_h_in_003_001-    1204858.1191073188
Rh003_008_001+    hidden_activ_out_h002_008    tia_h_in_003_001+    24777.472571937215
Rh003_008_001-    hidden_activ_out_h002_008    tia_h_in_003_001-    1195346.6123163868
Rh003_009_001+    hidden_activ_out_h002_009    tia_h_in_003_001+    30430.865871911952
Rh003_009_001-    hidden_activ_out_h002_009    tia_h_in_003_001-    1192665.9229089632
Rh003_010_001+    hidden_activ_out_h002_010    tia_h_in_003_001+    61559.2744377354
Rh003_010_001-    hidden_activ_out_h002_010    tia_h_in_003_001-    1205631.8939454013

* ----- Bias
    
        
Rb_h003_001+    b_003    tia_h_in_003_001+    1205714.7968574886
Rb_h003_001-    b_003    tia_h_in_003_001-    31045.31096155969


* ----- Difference (V(R+) - V(R-))

* Layer 000
* Neuron 1
Rh001_fb_001+     tia_h_in_001_001+ tia_h_out_001_001+ 6000
Rh001_fb_001-     tia_h_in_001_001- tia_h_out_001_001- 6000
XUh001_001+       0 tia_h_in_001_001+ Vcc+ Vcc- tia_h_out_001_001+ Ve OPA684_0
XUh001_001-       0 tia_h_in_001_001- Vcc+ Vcc- tia_h_out_001_001- Ve OPA684_0
Rh001_sum_001+    tia_h_out_001_001+ sum_h_in_001_001- 260
Rh001_sum_001-    tia_h_out_001_001- sum_h_in_001_001+ 260
Rh001_sum_l_001   sum_h_in_001_001+ 0 2020.9237114857817
Rh001_sum_fb_001  sum_h_in_001_001- sum_h_out_001_001 2020.9237114857817
XUh001_sum_001    sum_h_in_001_001+ sum_h_in_001_001- Vcc+ Vcc- sum_h_out_001_001 MAX4223
* Neuron 2
Rh001_fb_002+     tia_h_in_001_002+ tia_h_out_001_002+ 6000
Rh001_fb_002-     tia_h_in_001_002- tia_h_out_001_002- 6000
XUh001_002+       0 tia_h_in_001_002+ Vcc+ Vcc- tia_h_out_001_002+ Ve OPA684_0
XUh001_002-       0 tia_h_in_001_002- Vcc+ Vcc- tia_h_out_001_002- Ve OPA684_0
Rh001_sum_002+    tia_h_out_001_002+ sum_h_in_001_002- 260
Rh001_sum_002-    tia_h_out_001_002- sum_h_in_001_002+ 260
Rh001_sum_l_002   sum_h_in_001_002+ 0 2020.9237114857817
Rh001_sum_fb_002  sum_h_in_001_002- sum_h_out_001_002 2020.9237114857817
XUh001_sum_002    sum_h_in_001_002+ sum_h_in_001_002- Vcc+ Vcc- sum_h_out_001_002 MAX4223
* Neuron 3
Rh001_fb_003+     tia_h_in_001_003+ tia_h_out_001_003+ 6000
Rh001_fb_003-     tia_h_in_001_003- tia_h_out_001_003- 6000
XUh001_003+       0 tia_h_in_001_003+ Vcc+ Vcc- tia_h_out_001_003+ Ve OPA684_0
XUh001_003-       0 tia_h_in_001_003- Vcc+ Vcc- tia_h_out_001_003- Ve OPA684_0
Rh001_sum_003+    tia_h_out_001_003+ sum_h_in_001_003- 260
Rh001_sum_003-    tia_h_out_001_003- sum_h_in_001_003+ 260
Rh001_sum_l_003   sum_h_in_001_003+ 0 2020.9237114857817
Rh001_sum_fb_003  sum_h_in_001_003- sum_h_out_001_003 2020.9237114857817
XUh001_sum_003    sum_h_in_001_003+ sum_h_in_001_003- Vcc+ Vcc- sum_h_out_001_003 MAX4223
* Neuron 4
Rh001_fb_004+     tia_h_in_001_004+ tia_h_out_001_004+ 6000
Rh001_fb_004-     tia_h_in_001_004- tia_h_out_001_004- 6000
XUh001_004+       0 tia_h_in_001_004+ Vcc+ Vcc- tia_h_out_001_004+ Ve OPA684_0
XUh001_004-       0 tia_h_in_001_004- Vcc+ Vcc- tia_h_out_001_004- Ve OPA684_0
Rh001_sum_004+    tia_h_out_001_004+ sum_h_in_001_004- 260
Rh001_sum_004-    tia_h_out_001_004- sum_h_in_001_004+ 260
Rh001_sum_l_004   sum_h_in_001_004+ 0 2020.9237114857817
Rh001_sum_fb_004  sum_h_in_001_004- sum_h_out_001_004 2020.9237114857817
XUh001_sum_004    sum_h_in_001_004+ sum_h_in_001_004- Vcc+ Vcc- sum_h_out_001_004 MAX4223
* Neuron 5
Rh001_fb_005+     tia_h_in_001_005+ tia_h_out_001_005+ 6000
Rh001_fb_005-     tia_h_in_001_005- tia_h_out_001_005- 6000
XUh001_005+       0 tia_h_in_001_005+ Vcc+ Vcc- tia_h_out_001_005+ Ve OPA684_0
XUh001_005-       0 tia_h_in_001_005- Vcc+ Vcc- tia_h_out_001_005- Ve OPA684_0
Rh001_sum_005+    tia_h_out_001_005+ sum_h_in_001_005- 260
Rh001_sum_005-    tia_h_out_001_005- sum_h_in_001_005+ 260
Rh001_sum_l_005   sum_h_in_001_005+ 0 2020.9237114857817
Rh001_sum_fb_005  sum_h_in_001_005- sum_h_out_001_005 2020.9237114857817
XUh001_sum_005    sum_h_in_001_005+ sum_h_in_001_005- Vcc+ Vcc- sum_h_out_001_005 MAX4223
* Neuron 6
Rh001_fb_006+     tia_h_in_001_006+ tia_h_out_001_006+ 6000
Rh001_fb_006-     tia_h_in_001_006- tia_h_out_001_006- 6000
XUh001_006+       0 tia_h_in_001_006+ Vcc+ Vcc- tia_h_out_001_006+ Ve OPA684_0
XUh001_006-       0 tia_h_in_001_006- Vcc+ Vcc- tia_h_out_001_006- Ve OPA684_0
Rh001_sum_006+    tia_h_out_001_006+ sum_h_in_001_006- 260
Rh001_sum_006-    tia_h_out_001_006- sum_h_in_001_006+ 260
Rh001_sum_l_006   sum_h_in_001_006+ 0 2020.9237114857817
Rh001_sum_fb_006  sum_h_in_001_006- sum_h_out_001_006 2020.9237114857817
XUh001_sum_006    sum_h_in_001_006+ sum_h_in_001_006- Vcc+ Vcc- sum_h_out_001_006 MAX4223
* Neuron 7
Rh001_fb_007+     tia_h_in_001_007+ tia_h_out_001_007+ 6000
Rh001_fb_007-     tia_h_in_001_007- tia_h_out_001_007- 6000
XUh001_007+       0 tia_h_in_001_007+ Vcc+ Vcc- tia_h_out_001_007+ Ve OPA684_0
XUh001_007-       0 tia_h_in_001_007- Vcc+ Vcc- tia_h_out_001_007- Ve OPA684_0
Rh001_sum_007+    tia_h_out_001_007+ sum_h_in_001_007- 260
Rh001_sum_007-    tia_h_out_001_007- sum_h_in_001_007+ 260
Rh001_sum_l_007   sum_h_in_001_007+ 0 2020.9237114857817
Rh001_sum_fb_007  sum_h_in_001_007- sum_h_out_001_007 2020.9237114857817
XUh001_sum_007    sum_h_in_001_007+ sum_h_in_001_007- Vcc+ Vcc- sum_h_out_001_007 MAX4223
* Neuron 8
Rh001_fb_008+     tia_h_in_001_008+ tia_h_out_001_008+ 6000
Rh001_fb_008-     tia_h_in_001_008- tia_h_out_001_008- 6000
XUh001_008+       0 tia_h_in_001_008+ Vcc+ Vcc- tia_h_out_001_008+ Ve OPA684_0
XUh001_008-       0 tia_h_in_001_008- Vcc+ Vcc- tia_h_out_001_008- Ve OPA684_0
Rh001_sum_008+    tia_h_out_001_008+ sum_h_in_001_008- 260
Rh001_sum_008-    tia_h_out_001_008- sum_h_in_001_008+ 260
Rh001_sum_l_008   sum_h_in_001_008+ 0 2020.9237114857817
Rh001_sum_fb_008  sum_h_in_001_008- sum_h_out_001_008 2020.9237114857817
XUh001_sum_008    sum_h_in_001_008+ sum_h_in_001_008- Vcc+ Vcc- sum_h_out_001_008 MAX4223
* Neuron 9
Rh001_fb_009+     tia_h_in_001_009+ tia_h_out_001_009+ 6000
Rh001_fb_009-     tia_h_in_001_009- tia_h_out_001_009- 6000
XUh001_009+       0 tia_h_in_001_009+ Vcc+ Vcc- tia_h_out_001_009+ Ve OPA684_0
XUh001_009-       0 tia_h_in_001_009- Vcc+ Vcc- tia_h_out_001_009- Ve OPA684_0
Rh001_sum_009+    tia_h_out_001_009+ sum_h_in_001_009- 260
Rh001_sum_009-    tia_h_out_001_009- sum_h_in_001_009+ 260
Rh001_sum_l_009   sum_h_in_001_009+ 0 2020.9237114857817
Rh001_sum_fb_009  sum_h_in_001_009- sum_h_out_001_009 2020.9237114857817
XUh001_sum_009    sum_h_in_001_009+ sum_h_in_001_009- Vcc+ Vcc- sum_h_out_001_009 MAX4223
* Neuron 10
Rh001_fb_010+     tia_h_in_001_010+ tia_h_out_001_010+ 6000
Rh001_fb_010-     tia_h_in_001_010- tia_h_out_001_010- 6000
XUh001_010+       0 tia_h_in_001_010+ Vcc+ Vcc- tia_h_out_001_010+ Ve OPA684_0
XUh001_010-       0 tia_h_in_001_010- Vcc+ Vcc- tia_h_out_001_010- Ve OPA684_0
Rh001_sum_010+    tia_h_out_001_010+ sum_h_in_001_010- 260
Rh001_sum_010-    tia_h_out_001_010- sum_h_in_001_010+ 260
Rh001_sum_l_010   sum_h_in_001_010+ 0 2020.9237114857817
Rh001_sum_fb_010  sum_h_in_001_010- sum_h_out_001_010 2020.9237114857817
XUh001_sum_010    sum_h_in_001_010+ sum_h_in_001_010- Vcc+ Vcc- sum_h_out_001_010 MAX4223
* Neuron 11
Rh001_fb_011+     tia_h_in_001_011+ tia_h_out_001_011+ 6000
Rh001_fb_011-     tia_h_in_001_011- tia_h_out_001_011- 6000
XUh001_011+       0 tia_h_in_001_011+ Vcc+ Vcc- tia_h_out_001_011+ Ve OPA684_0
XUh001_011-       0 tia_h_in_001_011- Vcc+ Vcc- tia_h_out_001_011- Ve OPA684_0
Rh001_sum_011+    tia_h_out_001_011+ sum_h_in_001_011- 260
Rh001_sum_011-    tia_h_out_001_011- sum_h_in_001_011+ 260
Rh001_sum_l_011   sum_h_in_001_011+ 0 2020.9237114857817
Rh001_sum_fb_011  sum_h_in_001_011- sum_h_out_001_011 2020.9237114857817
XUh001_sum_011    sum_h_in_001_011+ sum_h_in_001_011- Vcc+ Vcc- sum_h_out_001_011 MAX4223
* Neuron 12
Rh001_fb_012+     tia_h_in_001_012+ tia_h_out_001_012+ 6000
Rh001_fb_012-     tia_h_in_001_012- tia_h_out_001_012- 6000
XUh001_012+       0 tia_h_in_001_012+ Vcc+ Vcc- tia_h_out_001_012+ Ve OPA684_0
XUh001_012-       0 tia_h_in_001_012- Vcc+ Vcc- tia_h_out_001_012- Ve OPA684_0
Rh001_sum_012+    tia_h_out_001_012+ sum_h_in_001_012- 260
Rh001_sum_012-    tia_h_out_001_012- sum_h_in_001_012+ 260
Rh001_sum_l_012   sum_h_in_001_012+ 0 2020.9237114857817
Rh001_sum_fb_012  sum_h_in_001_012- sum_h_out_001_012 2020.9237114857817
XUh001_sum_012    sum_h_in_001_012+ sum_h_in_001_012- Vcc+ Vcc- sum_h_out_001_012 MAX4223
* Neuron 13
Rh001_fb_013+     tia_h_in_001_013+ tia_h_out_001_013+ 6000
Rh001_fb_013-     tia_h_in_001_013- tia_h_out_001_013- 6000
XUh001_013+       0 tia_h_in_001_013+ Vcc+ Vcc- tia_h_out_001_013+ Ve OPA684_0
XUh001_013-       0 tia_h_in_001_013- Vcc+ Vcc- tia_h_out_001_013- Ve OPA684_0
Rh001_sum_013+    tia_h_out_001_013+ sum_h_in_001_013- 260
Rh001_sum_013-    tia_h_out_001_013- sum_h_in_001_013+ 260
Rh001_sum_l_013   sum_h_in_001_013+ 0 2020.9237114857817
Rh001_sum_fb_013  sum_h_in_001_013- sum_h_out_001_013 2020.9237114857817
XUh001_sum_013    sum_h_in_001_013+ sum_h_in_001_013- Vcc+ Vcc- sum_h_out_001_013 MAX4223
* Neuron 14
Rh001_fb_014+     tia_h_in_001_014+ tia_h_out_001_014+ 6000
Rh001_fb_014-     tia_h_in_001_014- tia_h_out_001_014- 6000
XUh001_014+       0 tia_h_in_001_014+ Vcc+ Vcc- tia_h_out_001_014+ Ve OPA684_0
XUh001_014-       0 tia_h_in_001_014- Vcc+ Vcc- tia_h_out_001_014- Ve OPA684_0
Rh001_sum_014+    tia_h_out_001_014+ sum_h_in_001_014- 260
Rh001_sum_014-    tia_h_out_001_014- sum_h_in_001_014+ 260
Rh001_sum_l_014   sum_h_in_001_014+ 0 2020.9237114857817
Rh001_sum_fb_014  sum_h_in_001_014- sum_h_out_001_014 2020.9237114857817
XUh001_sum_014    sum_h_in_001_014+ sum_h_in_001_014- Vcc+ Vcc- sum_h_out_001_014 MAX4223
* Neuron 15
Rh001_fb_015+     tia_h_in_001_015+ tia_h_out_001_015+ 6000
Rh001_fb_015-     tia_h_in_001_015- tia_h_out_001_015- 6000
XUh001_015+       0 tia_h_in_001_015+ Vcc+ Vcc- tia_h_out_001_015+ Ve OPA684_0
XUh001_015-       0 tia_h_in_001_015- Vcc+ Vcc- tia_h_out_001_015- Ve OPA684_0
Rh001_sum_015+    tia_h_out_001_015+ sum_h_in_001_015- 260
Rh001_sum_015-    tia_h_out_001_015- sum_h_in_001_015+ 260
Rh001_sum_l_015   sum_h_in_001_015+ 0 2020.9237114857817
Rh001_sum_fb_015  sum_h_in_001_015- sum_h_out_001_015 2020.9237114857817
XUh001_sum_015    sum_h_in_001_015+ sum_h_in_001_015- Vcc+ Vcc- sum_h_out_001_015 MAX4223
* Neuron 16
Rh001_fb_016+     tia_h_in_001_016+ tia_h_out_001_016+ 6000
Rh001_fb_016-     tia_h_in_001_016- tia_h_out_001_016- 6000
XUh001_016+       0 tia_h_in_001_016+ Vcc+ Vcc- tia_h_out_001_016+ Ve OPA684_0
XUh001_016-       0 tia_h_in_001_016- Vcc+ Vcc- tia_h_out_001_016- Ve OPA684_0
Rh001_sum_016+    tia_h_out_001_016+ sum_h_in_001_016- 260
Rh001_sum_016-    tia_h_out_001_016- sum_h_in_001_016+ 260
Rh001_sum_l_016   sum_h_in_001_016+ 0 2020.9237114857817
Rh001_sum_fb_016  sum_h_in_001_016- sum_h_out_001_016 2020.9237114857817
XUh001_sum_016    sum_h_in_001_016+ sum_h_in_001_016- Vcc+ Vcc- sum_h_out_001_016 MAX4223
* Neuron 17
Rh001_fb_017+     tia_h_in_001_017+ tia_h_out_001_017+ 6000
Rh001_fb_017-     tia_h_in_001_017- tia_h_out_001_017- 6000
XUh001_017+       0 tia_h_in_001_017+ Vcc+ Vcc- tia_h_out_001_017+ Ve OPA684_0
XUh001_017-       0 tia_h_in_001_017- Vcc+ Vcc- tia_h_out_001_017- Ve OPA684_0
Rh001_sum_017+    tia_h_out_001_017+ sum_h_in_001_017- 260
Rh001_sum_017-    tia_h_out_001_017- sum_h_in_001_017+ 260
Rh001_sum_l_017   sum_h_in_001_017+ 0 2020.9237114857817
Rh001_sum_fb_017  sum_h_in_001_017- sum_h_out_001_017 2020.9237114857817
XUh001_sum_017    sum_h_in_001_017+ sum_h_in_001_017- Vcc+ Vcc- sum_h_out_001_017 MAX4223
* Neuron 18
Rh001_fb_018+     tia_h_in_001_018+ tia_h_out_001_018+ 6000
Rh001_fb_018-     tia_h_in_001_018- tia_h_out_001_018- 6000
XUh001_018+       0 tia_h_in_001_018+ Vcc+ Vcc- tia_h_out_001_018+ Ve OPA684_0
XUh001_018-       0 tia_h_in_001_018- Vcc+ Vcc- tia_h_out_001_018- Ve OPA684_0
Rh001_sum_018+    tia_h_out_001_018+ sum_h_in_001_018- 260
Rh001_sum_018-    tia_h_out_001_018- sum_h_in_001_018+ 260
Rh001_sum_l_018   sum_h_in_001_018+ 0 2020.9237114857817
Rh001_sum_fb_018  sum_h_in_001_018- sum_h_out_001_018 2020.9237114857817
XUh001_sum_018    sum_h_in_001_018+ sum_h_in_001_018- Vcc+ Vcc- sum_h_out_001_018 MAX4223
* Neuron 19
Rh001_fb_019+     tia_h_in_001_019+ tia_h_out_001_019+ 6000
Rh001_fb_019-     tia_h_in_001_019- tia_h_out_001_019- 6000
XUh001_019+       0 tia_h_in_001_019+ Vcc+ Vcc- tia_h_out_001_019+ Ve OPA684_0
XUh001_019-       0 tia_h_in_001_019- Vcc+ Vcc- tia_h_out_001_019- Ve OPA684_0
Rh001_sum_019+    tia_h_out_001_019+ sum_h_in_001_019- 260
Rh001_sum_019-    tia_h_out_001_019- sum_h_in_001_019+ 260
Rh001_sum_l_019   sum_h_in_001_019+ 0 2020.9237114857817
Rh001_sum_fb_019  sum_h_in_001_019- sum_h_out_001_019 2020.9237114857817
XUh001_sum_019    sum_h_in_001_019+ sum_h_in_001_019- Vcc+ Vcc- sum_h_out_001_019 MAX4223
* Neuron 20
Rh001_fb_020+     tia_h_in_001_020+ tia_h_out_001_020+ 6000
Rh001_fb_020-     tia_h_in_001_020- tia_h_out_001_020- 6000
XUh001_020+       0 tia_h_in_001_020+ Vcc+ Vcc- tia_h_out_001_020+ Ve OPA684_0
XUh001_020-       0 tia_h_in_001_020- Vcc+ Vcc- tia_h_out_001_020- Ve OPA684_0
Rh001_sum_020+    tia_h_out_001_020+ sum_h_in_001_020- 260
Rh001_sum_020-    tia_h_out_001_020- sum_h_in_001_020+ 260
Rh001_sum_l_020   sum_h_in_001_020+ 0 2020.9237114857817
Rh001_sum_fb_020  sum_h_in_001_020- sum_h_out_001_020 2020.9237114857817
XUh001_sum_020    sum_h_in_001_020+ sum_h_in_001_020- Vcc+ Vcc- sum_h_out_001_020 MAX4223

* Layer 001
* Neuron 1
Rh002_fb_001+     tia_h_in_002_001+ tia_h_out_002_001+ 6000
Rh002_fb_001-     tia_h_in_002_001- tia_h_out_002_001- 6000
XUh002_001+       0 tia_h_in_002_001+ Vcc+ Vcc- tia_h_out_002_001+ Ve OPA684_0
XUh002_001-       0 tia_h_in_002_001- Vcc+ Vcc- tia_h_out_002_001- Ve OPA684_0
Rh002_sum_001+    tia_h_out_002_001+ sum_h_in_002_001- 260
Rh002_sum_001-    tia_h_out_002_001- sum_h_in_002_001+ 260
Rh002_sum_l_001   sum_h_in_002_001+ 0 2020.9237114857817
Rh002_sum_fb_001  sum_h_in_002_001- sum_h_out_002_001 2020.9237114857817
XUh002_sum_001    sum_h_in_002_001+ sum_h_in_002_001- Vcc+ Vcc- sum_h_out_002_001 MAX4223
* Neuron 2
Rh002_fb_002+     tia_h_in_002_002+ tia_h_out_002_002+ 6000
Rh002_fb_002-     tia_h_in_002_002- tia_h_out_002_002- 6000
XUh002_002+       0 tia_h_in_002_002+ Vcc+ Vcc- tia_h_out_002_002+ Ve OPA684_0
XUh002_002-       0 tia_h_in_002_002- Vcc+ Vcc- tia_h_out_002_002- Ve OPA684_0
Rh002_sum_002+    tia_h_out_002_002+ sum_h_in_002_002- 260
Rh002_sum_002-    tia_h_out_002_002- sum_h_in_002_002+ 260
Rh002_sum_l_002   sum_h_in_002_002+ 0 2020.9237114857817
Rh002_sum_fb_002  sum_h_in_002_002- sum_h_out_002_002 2020.9237114857817
XUh002_sum_002    sum_h_in_002_002+ sum_h_in_002_002- Vcc+ Vcc- sum_h_out_002_002 MAX4223
* Neuron 3
Rh002_fb_003+     tia_h_in_002_003+ tia_h_out_002_003+ 6000
Rh002_fb_003-     tia_h_in_002_003- tia_h_out_002_003- 6000
XUh002_003+       0 tia_h_in_002_003+ Vcc+ Vcc- tia_h_out_002_003+ Ve OPA684_0
XUh002_003-       0 tia_h_in_002_003- Vcc+ Vcc- tia_h_out_002_003- Ve OPA684_0
Rh002_sum_003+    tia_h_out_002_003+ sum_h_in_002_003- 260
Rh002_sum_003-    tia_h_out_002_003- sum_h_in_002_003+ 260
Rh002_sum_l_003   sum_h_in_002_003+ 0 2020.9237114857817
Rh002_sum_fb_003  sum_h_in_002_003- sum_h_out_002_003 2020.9237114857817
XUh002_sum_003    sum_h_in_002_003+ sum_h_in_002_003- Vcc+ Vcc- sum_h_out_002_003 MAX4223
* Neuron 4
Rh002_fb_004+     tia_h_in_002_004+ tia_h_out_002_004+ 6000
Rh002_fb_004-     tia_h_in_002_004- tia_h_out_002_004- 6000
XUh002_004+       0 tia_h_in_002_004+ Vcc+ Vcc- tia_h_out_002_004+ Ve OPA684_0
XUh002_004-       0 tia_h_in_002_004- Vcc+ Vcc- tia_h_out_002_004- Ve OPA684_0
Rh002_sum_004+    tia_h_out_002_004+ sum_h_in_002_004- 260
Rh002_sum_004-    tia_h_out_002_004- sum_h_in_002_004+ 260
Rh002_sum_l_004   sum_h_in_002_004+ 0 2020.9237114857817
Rh002_sum_fb_004  sum_h_in_002_004- sum_h_out_002_004 2020.9237114857817
XUh002_sum_004    sum_h_in_002_004+ sum_h_in_002_004- Vcc+ Vcc- sum_h_out_002_004 MAX4223
* Neuron 5
Rh002_fb_005+     tia_h_in_002_005+ tia_h_out_002_005+ 6000
Rh002_fb_005-     tia_h_in_002_005- tia_h_out_002_005- 6000
XUh002_005+       0 tia_h_in_002_005+ Vcc+ Vcc- tia_h_out_002_005+ Ve OPA684_0
XUh002_005-       0 tia_h_in_002_005- Vcc+ Vcc- tia_h_out_002_005- Ve OPA684_0
Rh002_sum_005+    tia_h_out_002_005+ sum_h_in_002_005- 260
Rh002_sum_005-    tia_h_out_002_005- sum_h_in_002_005+ 260
Rh002_sum_l_005   sum_h_in_002_005+ 0 2020.9237114857817
Rh002_sum_fb_005  sum_h_in_002_005- sum_h_out_002_005 2020.9237114857817
XUh002_sum_005    sum_h_in_002_005+ sum_h_in_002_005- Vcc+ Vcc- sum_h_out_002_005 MAX4223
* Neuron 6
Rh002_fb_006+     tia_h_in_002_006+ tia_h_out_002_006+ 6000
Rh002_fb_006-     tia_h_in_002_006- tia_h_out_002_006- 6000
XUh002_006+       0 tia_h_in_002_006+ Vcc+ Vcc- tia_h_out_002_006+ Ve OPA684_0
XUh002_006-       0 tia_h_in_002_006- Vcc+ Vcc- tia_h_out_002_006- Ve OPA684_0
Rh002_sum_006+    tia_h_out_002_006+ sum_h_in_002_006- 260
Rh002_sum_006-    tia_h_out_002_006- sum_h_in_002_006+ 260
Rh002_sum_l_006   sum_h_in_002_006+ 0 2020.9237114857817
Rh002_sum_fb_006  sum_h_in_002_006- sum_h_out_002_006 2020.9237114857817
XUh002_sum_006    sum_h_in_002_006+ sum_h_in_002_006- Vcc+ Vcc- sum_h_out_002_006 MAX4223
* Neuron 7
Rh002_fb_007+     tia_h_in_002_007+ tia_h_out_002_007+ 6000
Rh002_fb_007-     tia_h_in_002_007- tia_h_out_002_007- 6000
XUh002_007+       0 tia_h_in_002_007+ Vcc+ Vcc- tia_h_out_002_007+ Ve OPA684_0
XUh002_007-       0 tia_h_in_002_007- Vcc+ Vcc- tia_h_out_002_007- Ve OPA684_0
Rh002_sum_007+    tia_h_out_002_007+ sum_h_in_002_007- 260
Rh002_sum_007-    tia_h_out_002_007- sum_h_in_002_007+ 260
Rh002_sum_l_007   sum_h_in_002_007+ 0 2020.9237114857817
Rh002_sum_fb_007  sum_h_in_002_007- sum_h_out_002_007 2020.9237114857817
XUh002_sum_007    sum_h_in_002_007+ sum_h_in_002_007- Vcc+ Vcc- sum_h_out_002_007 MAX4223
* Neuron 8
Rh002_fb_008+     tia_h_in_002_008+ tia_h_out_002_008+ 6000
Rh002_fb_008-     tia_h_in_002_008- tia_h_out_002_008- 6000
XUh002_008+       0 tia_h_in_002_008+ Vcc+ Vcc- tia_h_out_002_008+ Ve OPA684_0
XUh002_008-       0 tia_h_in_002_008- Vcc+ Vcc- tia_h_out_002_008- Ve OPA684_0
Rh002_sum_008+    tia_h_out_002_008+ sum_h_in_002_008- 260
Rh002_sum_008-    tia_h_out_002_008- sum_h_in_002_008+ 260
Rh002_sum_l_008   sum_h_in_002_008+ 0 2020.9237114857817
Rh002_sum_fb_008  sum_h_in_002_008- sum_h_out_002_008 2020.9237114857817
XUh002_sum_008    sum_h_in_002_008+ sum_h_in_002_008- Vcc+ Vcc- sum_h_out_002_008 MAX4223
* Neuron 9
Rh002_fb_009+     tia_h_in_002_009+ tia_h_out_002_009+ 6000
Rh002_fb_009-     tia_h_in_002_009- tia_h_out_002_009- 6000
XUh002_009+       0 tia_h_in_002_009+ Vcc+ Vcc- tia_h_out_002_009+ Ve OPA684_0
XUh002_009-       0 tia_h_in_002_009- Vcc+ Vcc- tia_h_out_002_009- Ve OPA684_0
Rh002_sum_009+    tia_h_out_002_009+ sum_h_in_002_009- 260
Rh002_sum_009-    tia_h_out_002_009- sum_h_in_002_009+ 260
Rh002_sum_l_009   sum_h_in_002_009+ 0 2020.9237114857817
Rh002_sum_fb_009  sum_h_in_002_009- sum_h_out_002_009 2020.9237114857817
XUh002_sum_009    sum_h_in_002_009+ sum_h_in_002_009- Vcc+ Vcc- sum_h_out_002_009 MAX4223
* Neuron 10
Rh002_fb_010+     tia_h_in_002_010+ tia_h_out_002_010+ 6000
Rh002_fb_010-     tia_h_in_002_010- tia_h_out_002_010- 6000
XUh002_010+       0 tia_h_in_002_010+ Vcc+ Vcc- tia_h_out_002_010+ Ve OPA684_0
XUh002_010-       0 tia_h_in_002_010- Vcc+ Vcc- tia_h_out_002_010- Ve OPA684_0
Rh002_sum_010+    tia_h_out_002_010+ sum_h_in_002_010- 260
Rh002_sum_010-    tia_h_out_002_010- sum_h_in_002_010+ 260
Rh002_sum_l_010   sum_h_in_002_010+ 0 2020.9237114857817
Rh002_sum_fb_010  sum_h_in_002_010- sum_h_out_002_010 2020.9237114857817
XUh002_sum_010    sum_h_in_002_010+ sum_h_in_002_010- Vcc+ Vcc- sum_h_out_002_010 MAX4223

* Layer 002
* Neuron 1
Rh003_fb_001+     tia_h_in_003_001+ tia_h_out_003_001+ 6000
Rh003_fb_001-     tia_h_in_003_001- tia_h_out_003_001- 6000
XUh003_001+       0 tia_h_in_003_001+ Vcc+ Vcc- tia_h_out_003_001+ Ve OPA684_0
XUh003_001-       0 tia_h_in_003_001- Vcc+ Vcc- tia_h_out_003_001- Ve OPA684_0
Rh003_sum_001+    tia_h_out_003_001+ sum_h_in_003_001- 260
Rh003_sum_001-    tia_h_out_003_001- sum_h_in_003_001+ 260
Rh003_sum_l_001   sum_h_in_003_001+ 0 2020.9237114857817
Rh003_sum_fb_001  sum_h_in_003_001- sum_h_out_003_001 2020.9237114857817
XUh003_sum_001    sum_h_in_003_001+ sum_h_in_003_001- Vcc+ Vcc- sum_h_out_003_001 MAX4223


* ----- Activation function Hard-Tanh)


* Layer 000
* Neuron 1
* XHardTanh_h001_001 sum_h_out_001_001 hidden_activ_out_h001_001 HardTanh PARAMS: V_clip=-0.3
XReLU_001_001 sum_h_out_001_001 hidden_activ_out_h001_001 ReLU
*XSigmoid_001_001 sum_h_out_001_001 hidden_activ_out_h001_001 RNN_Sigmoid3_HA
* Neuron 2
* XHardTanh_h001_002 sum_h_out_001_002 hidden_activ_out_h001_002 HardTanh PARAMS: V_clip=-0.3
XReLU_001_002 sum_h_out_001_002 hidden_activ_out_h001_002 ReLU
*XSigmoid_001_002 sum_h_out_001_002 hidden_activ_out_h001_002 RNN_Sigmoid3_HA
* Neuron 3
* XHardTanh_h001_003 sum_h_out_001_003 hidden_activ_out_h001_003 HardTanh PARAMS: V_clip=-0.3
XReLU_001_003 sum_h_out_001_003 hidden_activ_out_h001_003 ReLU
*XSigmoid_001_003 sum_h_out_001_003 hidden_activ_out_h001_003 RNN_Sigmoid3_HA
* Neuron 4
* XHardTanh_h001_004 sum_h_out_001_004 hidden_activ_out_h001_004 HardTanh PARAMS: V_clip=-0.3
XReLU_001_004 sum_h_out_001_004 hidden_activ_out_h001_004 ReLU
*XSigmoid_001_004 sum_h_out_001_004 hidden_activ_out_h001_004 RNN_Sigmoid3_HA
* Neuron 5
* XHardTanh_h001_005 sum_h_out_001_005 hidden_activ_out_h001_005 HardTanh PARAMS: V_clip=-0.3
XReLU_001_005 sum_h_out_001_005 hidden_activ_out_h001_005 ReLU
*XSigmoid_001_005 sum_h_out_001_005 hidden_activ_out_h001_005 RNN_Sigmoid3_HA
* Neuron 6
* XHardTanh_h001_006 sum_h_out_001_006 hidden_activ_out_h001_006 HardTanh PARAMS: V_clip=-0.3
XReLU_001_006 sum_h_out_001_006 hidden_activ_out_h001_006 ReLU
*XSigmoid_001_006 sum_h_out_001_006 hidden_activ_out_h001_006 RNN_Sigmoid3_HA
* Neuron 7
* XHardTanh_h001_007 sum_h_out_001_007 hidden_activ_out_h001_007 HardTanh PARAMS: V_clip=-0.3
XReLU_001_007 sum_h_out_001_007 hidden_activ_out_h001_007 ReLU
*XSigmoid_001_007 sum_h_out_001_007 hidden_activ_out_h001_007 RNN_Sigmoid3_HA
* Neuron 8
* XHardTanh_h001_008 sum_h_out_001_008 hidden_activ_out_h001_008 HardTanh PARAMS: V_clip=-0.3
XReLU_001_008 sum_h_out_001_008 hidden_activ_out_h001_008 ReLU
*XSigmoid_001_008 sum_h_out_001_008 hidden_activ_out_h001_008 RNN_Sigmoid3_HA
* Neuron 9
* XHardTanh_h001_009 sum_h_out_001_009 hidden_activ_out_h001_009 HardTanh PARAMS: V_clip=-0.3
XReLU_001_009 sum_h_out_001_009 hidden_activ_out_h001_009 ReLU
*XSigmoid_001_009 sum_h_out_001_009 hidden_activ_out_h001_009 RNN_Sigmoid3_HA
* Neuron 10
* XHardTanh_h001_010 sum_h_out_001_010 hidden_activ_out_h001_010 HardTanh PARAMS: V_clip=-0.3
XReLU_001_010 sum_h_out_001_010 hidden_activ_out_h001_010 ReLU
*XSigmoid_001_010 sum_h_out_001_010 hidden_activ_out_h001_010 RNN_Sigmoid3_HA
* Neuron 11
* XHardTanh_h001_011 sum_h_out_001_011 hidden_activ_out_h001_011 HardTanh PARAMS: V_clip=-0.3
XReLU_001_011 sum_h_out_001_011 hidden_activ_out_h001_011 ReLU
*XSigmoid_001_011 sum_h_out_001_011 hidden_activ_out_h001_011 RNN_Sigmoid3_HA
* Neuron 12
* XHardTanh_h001_012 sum_h_out_001_012 hidden_activ_out_h001_012 HardTanh PARAMS: V_clip=-0.3
XReLU_001_012 sum_h_out_001_012 hidden_activ_out_h001_012 ReLU
*XSigmoid_001_012 sum_h_out_001_012 hidden_activ_out_h001_012 RNN_Sigmoid3_HA
* Neuron 13
* XHardTanh_h001_013 sum_h_out_001_013 hidden_activ_out_h001_013 HardTanh PARAMS: V_clip=-0.3
XReLU_001_013 sum_h_out_001_013 hidden_activ_out_h001_013 ReLU
*XSigmoid_001_013 sum_h_out_001_013 hidden_activ_out_h001_013 RNN_Sigmoid3_HA
* Neuron 14
* XHardTanh_h001_014 sum_h_out_001_014 hidden_activ_out_h001_014 HardTanh PARAMS: V_clip=-0.3
XReLU_001_014 sum_h_out_001_014 hidden_activ_out_h001_014 ReLU
*XSigmoid_001_014 sum_h_out_001_014 hidden_activ_out_h001_014 RNN_Sigmoid3_HA
* Neuron 15
* XHardTanh_h001_015 sum_h_out_001_015 hidden_activ_out_h001_015 HardTanh PARAMS: V_clip=-0.3
XReLU_001_015 sum_h_out_001_015 hidden_activ_out_h001_015 ReLU
*XSigmoid_001_015 sum_h_out_001_015 hidden_activ_out_h001_015 RNN_Sigmoid3_HA
* Neuron 16
* XHardTanh_h001_016 sum_h_out_001_016 hidden_activ_out_h001_016 HardTanh PARAMS: V_clip=-0.3
XReLU_001_016 sum_h_out_001_016 hidden_activ_out_h001_016 ReLU
*XSigmoid_001_016 sum_h_out_001_016 hidden_activ_out_h001_016 RNN_Sigmoid3_HA
* Neuron 17
* XHardTanh_h001_017 sum_h_out_001_017 hidden_activ_out_h001_017 HardTanh PARAMS: V_clip=-0.3
XReLU_001_017 sum_h_out_001_017 hidden_activ_out_h001_017 ReLU
*XSigmoid_001_017 sum_h_out_001_017 hidden_activ_out_h001_017 RNN_Sigmoid3_HA
* Neuron 18
* XHardTanh_h001_018 sum_h_out_001_018 hidden_activ_out_h001_018 HardTanh PARAMS: V_clip=-0.3
XReLU_001_018 sum_h_out_001_018 hidden_activ_out_h001_018 ReLU
*XSigmoid_001_018 sum_h_out_001_018 hidden_activ_out_h001_018 RNN_Sigmoid3_HA
* Neuron 19
* XHardTanh_h001_019 sum_h_out_001_019 hidden_activ_out_h001_019 HardTanh PARAMS: V_clip=-0.3
XReLU_001_019 sum_h_out_001_019 hidden_activ_out_h001_019 ReLU
*XSigmoid_001_019 sum_h_out_001_019 hidden_activ_out_h001_019 RNN_Sigmoid3_HA
* Neuron 20
* XHardTanh_h001_020 sum_h_out_001_020 hidden_activ_out_h001_020 HardTanh PARAMS: V_clip=-0.3
XReLU_001_020 sum_h_out_001_020 hidden_activ_out_h001_020 ReLU
*XSigmoid_001_020 sum_h_out_001_020 hidden_activ_out_h001_020 RNN_Sigmoid3_HA

* Layer 001
* Neuron 1
* XHardTanh_h002_001 sum_h_out_002_001 hidden_activ_out_h002_001 HardTanh PARAMS: V_clip=-0.3
XReLU_002_001 sum_h_out_002_001 hidden_activ_out_h002_001 ReLU
*XSigmoid_002_001 sum_h_out_002_001 hidden_activ_out_h002_001 RNN_Sigmoid3_HA
* Neuron 2
* XHardTanh_h002_002 sum_h_out_002_002 hidden_activ_out_h002_002 HardTanh PARAMS: V_clip=-0.3
XReLU_002_002 sum_h_out_002_002 hidden_activ_out_h002_002 ReLU
*XSigmoid_002_002 sum_h_out_002_002 hidden_activ_out_h002_002 RNN_Sigmoid3_HA
* Neuron 3
* XHardTanh_h002_003 sum_h_out_002_003 hidden_activ_out_h002_003 HardTanh PARAMS: V_clip=-0.3
XReLU_002_003 sum_h_out_002_003 hidden_activ_out_h002_003 ReLU
*XSigmoid_002_003 sum_h_out_002_003 hidden_activ_out_h002_003 RNN_Sigmoid3_HA
* Neuron 4
* XHardTanh_h002_004 sum_h_out_002_004 hidden_activ_out_h002_004 HardTanh PARAMS: V_clip=-0.3
XReLU_002_004 sum_h_out_002_004 hidden_activ_out_h002_004 ReLU
*XSigmoid_002_004 sum_h_out_002_004 hidden_activ_out_h002_004 RNN_Sigmoid3_HA
* Neuron 5
* XHardTanh_h002_005 sum_h_out_002_005 hidden_activ_out_h002_005 HardTanh PARAMS: V_clip=-0.3
XReLU_002_005 sum_h_out_002_005 hidden_activ_out_h002_005 ReLU
*XSigmoid_002_005 sum_h_out_002_005 hidden_activ_out_h002_005 RNN_Sigmoid3_HA
* Neuron 6
* XHardTanh_h002_006 sum_h_out_002_006 hidden_activ_out_h002_006 HardTanh PARAMS: V_clip=-0.3
XReLU_002_006 sum_h_out_002_006 hidden_activ_out_h002_006 ReLU
*XSigmoid_002_006 sum_h_out_002_006 hidden_activ_out_h002_006 RNN_Sigmoid3_HA
* Neuron 7
* XHardTanh_h002_007 sum_h_out_002_007 hidden_activ_out_h002_007 HardTanh PARAMS: V_clip=-0.3
XReLU_002_007 sum_h_out_002_007 hidden_activ_out_h002_007 ReLU
*XSigmoid_002_007 sum_h_out_002_007 hidden_activ_out_h002_007 RNN_Sigmoid3_HA
* Neuron 8
* XHardTanh_h002_008 sum_h_out_002_008 hidden_activ_out_h002_008 HardTanh PARAMS: V_clip=-0.3
XReLU_002_008 sum_h_out_002_008 hidden_activ_out_h002_008 ReLU
*XSigmoid_002_008 sum_h_out_002_008 hidden_activ_out_h002_008 RNN_Sigmoid3_HA
* Neuron 9
* XHardTanh_h002_009 sum_h_out_002_009 hidden_activ_out_h002_009 HardTanh PARAMS: V_clip=-0.3
XReLU_002_009 sum_h_out_002_009 hidden_activ_out_h002_009 ReLU
*XSigmoid_002_009 sum_h_out_002_009 hidden_activ_out_h002_009 RNN_Sigmoid3_HA
* Neuron 10
* XHardTanh_h002_010 sum_h_out_002_010 hidden_activ_out_h002_010 HardTanh PARAMS: V_clip=-0.3
XReLU_002_010 sum_h_out_002_010 hidden_activ_out_h002_010 ReLU
*XSigmoid_002_010 sum_h_out_002_010 hidden_activ_out_h002_010 RNN_Sigmoid3_HA

* Layer 002
* Neuron 1
* XHardTanh_h003_001 sum_h_out_003_001 hidden_activ_out_h003_001 HardTanh PARAMS: V_clip=-0.3
XReLU_003_001 sum_h_out_003_001 hidden_activ_out_h003_001 ReLU
*XSigmoid_003_001 sum_h_out_003_001 hidden_activ_out_h003_001 RNN_Sigmoid3_HA


.END