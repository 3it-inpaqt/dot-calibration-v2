* Netlist that describe the physical circuit (components and connexions between them) to simulate, in Xyce formalism.
* To make the translation from any network size, the circuit is scaled up automatically using Jinja template engine.
*
* Xyce: https://xyce.sandia.gov
* Jinja: https://jinja.palletsprojects.com

* ======================== Simulation parameters ==========================
.param simtime=420n
.TRAN 0.20ns {simtime}

* OPTIONS TIMEINT change the time integration parameters
* ERROPTION (If 0 Local Truncation Error is used)
* METHOD: Time integration method
* NLMIN, NLMAX:  lower and upper bound for the desired number of nonlinear iterations
* DELMAX: The maximum time step-size used
* This additional line allows to fix convergence problem but increases the simulation time
*.OPTIONS TIMEINT ERROPTION=1 METHOD=GEAR NLMIN=3 NLMAX=8 DELMAX=1.0e-10
*.OPTIONS ERROPTION=1 METHOD=GEAR NLMIN=3 NLMAX=8 DELMAX=1.0e-10

* List variables to save in the result table
.PRINT TRAN V(sum_h_out_002_001) V(hidden_activ_out_h002_001)
+ V(i_001) V(i_002) V(i_003) V(i_004) V(i_005) V(i_006) V(i_007) V(i_008) V(i_009) V(i_010) V(i_011) V(i_012) V(i_013) V(i_014) V(i_015) V(i_016) V(i_017) V(i_018) V(i_019) V(i_020) V(i_021) V(i_022) V(i_023) V(i_024) V(i_025)
+ V(sum_h_out_001_001) V(hidden_activ_out_h001_001) V(sum_h_out_001_002) V(hidden_activ_out_h001_002) V(sum_h_out_001_003) V(hidden_activ_out_h001_003) V(sum_h_out_001_004) V(hidden_activ_out_h001_004) V(sum_h_out_001_005) V(hidden_activ_out_h001_005)
+ V(tia_h_out_001_001+) V(tia_h_out_001_001-) V(tia_h_out_001_002+) V(tia_h_out_001_002-) V(tia_h_out_001_003+) V(tia_h_out_001_003-) V(tia_h_out_001_004+) V(tia_h_out_001_004-) V(tia_h_out_001_005+) V(tia_h_out_001_005-)
+ V(b_001)
+ V(sum_h_out_002_001) V(hidden_activ_out_h002_001)
+ V(tia_h_out_002_001+) V(tia_h_out_002_001-)
+ V(b_002)

* =============================== Models ==================================

* Call the defined components model from the specified path
*.INCLUDE "./components/MAX4223.sub"
.INCLUDE "./components/TLV3501.sub"
*.INCLUDE "./components/OPA684.sub"

* Import custom sub-circuits
.INCLUDE "./components/activations.sub"
.INCLUDE "./components/lumped_line.sub"

* Define diode model
.MODEL D_BAV74_1 D( IS=2.073F N=1 BV=50 IBV=100N RS=1.336
+      CJO=2P VJ=750M M=330M FC=500M TT=5.771N
+      EG=1.11 XTI=3 KF=0 AF=1 )

* ============================== Voltages =================================

* ----- Input pulses
* Vi_num: The input voltage as pulse sequences
Vi_001    i_001    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_002    i_002    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_003    i_003    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_004    i_004    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_005    i_005    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_006    i_006    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_007    i_007    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_008    i_008    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_009    i_009    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_010    i_010    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_011    i_011    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_012    i_012    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_013    i_013    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_014    i_014    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_015    i_015    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_016    i_016    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_017    i_017    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_018    i_018    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_019    i_019    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_020    i_020    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_021    i_021    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_022    i_022    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_023    i_023    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.200V 400.00ns 0.200V 401.00ns 0.000V
Vi_024    i_024    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V
Vi_025    i_025    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.000V 400.00ns 0.000V 401.00ns 0.000V

* Vb_num: The bias voltage as pulse sequences

Vb_001    b_001    0    PWL 0.00ns 0.000V 1.00ns 0.000V 2.00ns 0.200V 400.00ns 0.200V 401.00ns 0.000V
Vb_002    b_002    0    PWL 0.00ns 0.000V 11.00ns 0.000V 12.00ns 0.200V 410.00ns 0.200V 411.00ns 0.000V

Ve        Ve       0    3
Vcc-      Vcc-     0    -5
Vcc+      Vcc+     0    5

* ============================ NN Parameters ==============================
* Parameters (weights and bias) naming convention: "Rl_i_j+" where:
*   R: Always "R" to inform Xyce it is a resistance
*   l: layer name, "h" for the hidden and output layers and "b" for the biases.
*   i: index of the weight of a neuron (start from 1)
*   j: index of the neuron (start from 1)
*   +: parameter polarity, + or -

* ----------------------------- Layers -----------------------------


* ----- Weights
* Layer 001

* Neuron 1
Rh001_001_001+    i_001    tia_h_in_001_001+    15000
Rh001_001_001-    i_001    tia_h_in_001_001-    12488
Rh001_002_001+    i_002    tia_h_in_001_001+    15000
Rh001_002_001-    i_002    tia_h_in_001_001-    10890
Rh001_003_001+    i_003    tia_h_in_001_001+    15000
Rh001_003_001-    i_003    tia_h_in_001_001-    10897
Rh001_004_001+    i_004    tia_h_in_001_001+    15000
Rh001_004_001-    i_004    tia_h_in_001_001-    13122
Rh001_005_001+    i_005    tia_h_in_001_001+    15000
Rh001_005_001-    i_005    tia_h_in_001_001-    13804
Rh001_006_001+    i_006    tia_h_in_001_001+    15000
Rh001_006_001-    i_006    tia_h_in_001_001-    13176
Rh001_007_001+    i_007    tia_h_in_001_001+    15000
Rh001_007_001-    i_007    tia_h_in_001_001-    14611
Rh001_008_001+    i_008    tia_h_in_001_001+    15000
Rh001_008_001-    i_008    tia_h_in_001_001-    13908
Rh001_009_001+    i_009    tia_h_in_001_001+    15000
Rh001_009_001-    i_009    tia_h_in_001_001-    13680
Rh001_010_001+    i_010    tia_h_in_001_001+    15000
Rh001_010_001-    i_010    tia_h_in_001_001-    12903
Rh001_011_001+    i_011    tia_h_in_001_001+    15000
Rh001_011_001-    i_011    tia_h_in_001_001-    11045
Rh001_012_001+    i_012    tia_h_in_001_001+    15000
Rh001_012_001-    i_012    tia_h_in_001_001-    12559
Rh001_013_001+    i_013    tia_h_in_001_001+    15000
Rh001_013_001-    i_013    tia_h_in_001_001-    14041
Rh001_014_001+    i_014    tia_h_in_001_001+    15000
Rh001_014_001-    i_014    tia_h_in_001_001-    12246
Rh001_015_001+    i_015    tia_h_in_001_001+    15000
Rh001_015_001-    i_015    tia_h_in_001_001-    11312
Rh001_016_001+    i_016    tia_h_in_001_001+    15000
Rh001_016_001-    i_016    tia_h_in_001_001-    12751
Rh001_017_001+    i_017    tia_h_in_001_001+    15000
Rh001_017_001-    i_017    tia_h_in_001_001-    11724
Rh001_018_001+    i_018    tia_h_in_001_001+    15000
Rh001_018_001-    i_018    tia_h_in_001_001-    11368
Rh001_019_001+    i_019    tia_h_in_001_001+    15000
Rh001_019_001-    i_019    tia_h_in_001_001-    12228
Rh001_020_001+    i_020    tia_h_in_001_001+    15000
Rh001_020_001-    i_020    tia_h_in_001_001-    12546
Rh001_021_001+    i_021    tia_h_in_001_001+    15000
Rh001_021_001-    i_021    tia_h_in_001_001-    11168
Rh001_022_001+    i_022    tia_h_in_001_001+    15000
Rh001_022_001-    i_022    tia_h_in_001_001-    11641
Rh001_023_001+    i_023    tia_h_in_001_001+    15000
Rh001_023_001-    i_023    tia_h_in_001_001-    12108
Rh001_024_001+    i_024    tia_h_in_001_001+    15000
Rh001_024_001-    i_024    tia_h_in_001_001-    11903
Rh001_025_001+    i_025    tia_h_in_001_001+    15000
Rh001_025_001-    i_025    tia_h_in_001_001-    12139

* Neuron 2
Rh001_001_002+    i_001    tia_h_in_001_002+    15000
Rh001_001_002-    i_001    tia_h_in_001_002-    9078
Rh001_002_002+    i_002    tia_h_in_001_002+    15000
Rh001_002_002-    i_002    tia_h_in_001_002-    9589
Rh001_003_002+    i_003    tia_h_in_001_002+    15000
Rh001_003_002-    i_003    tia_h_in_001_002-    9539
Rh001_004_002+    i_004    tia_h_in_001_002+    15000
Rh001_004_002-    i_004    tia_h_in_001_002-    9676
Rh001_005_002+    i_005    tia_h_in_001_002+    15000
Rh001_005_002-    i_005    tia_h_in_001_002-    9301
Rh001_006_002+    i_006    tia_h_in_001_002+    15000
Rh001_006_002-    i_006    tia_h_in_001_002-    9436
Rh001_007_002+    i_007    tia_h_in_001_002+    15000
Rh001_007_002-    i_007    tia_h_in_001_002-    9505
Rh001_008_002+    i_008    tia_h_in_001_002+    15000
Rh001_008_002-    i_008    tia_h_in_001_002-    9602
Rh001_009_002+    i_009    tia_h_in_001_002+    15000
Rh001_009_002-    i_009    tia_h_in_001_002-    10011
Rh001_010_002+    i_010    tia_h_in_001_002+    15000
Rh001_010_002-    i_010    tia_h_in_001_002-    9476
Rh001_011_002+    i_011    tia_h_in_001_002+    15000
Rh001_011_002-    i_011    tia_h_in_001_002-    9372
Rh001_012_002+    i_012    tia_h_in_001_002+    15000
Rh001_012_002-    i_012    tia_h_in_001_002-    9462
Rh001_013_002+    i_013    tia_h_in_001_002+    15000
Rh001_013_002-    i_013    tia_h_in_001_002-    9497
Rh001_014_002+    i_014    tia_h_in_001_002+    15000
Rh001_014_002-    i_014    tia_h_in_001_002-    9618
Rh001_015_002+    i_015    tia_h_in_001_002+    15000
Rh001_015_002-    i_015    tia_h_in_001_002-    9797
Rh001_016_002+    i_016    tia_h_in_001_002+    15000
Rh001_016_002-    i_016    tia_h_in_001_002-    9665
Rh001_017_002+    i_017    tia_h_in_001_002+    15000
Rh001_017_002-    i_017    tia_h_in_001_002-    9408
Rh001_018_002+    i_018    tia_h_in_001_002+    15000
Rh001_018_002-    i_018    tia_h_in_001_002-    9533
Rh001_019_002+    i_019    tia_h_in_001_002+    15000
Rh001_019_002-    i_019    tia_h_in_001_002-    9452
Rh001_020_002+    i_020    tia_h_in_001_002+    15000
Rh001_020_002-    i_020    tia_h_in_001_002-    9352
Rh001_021_002+    i_021    tia_h_in_001_002+    15000
Rh001_021_002-    i_021    tia_h_in_001_002-    9297
Rh001_022_002+    i_022    tia_h_in_001_002+    15000
Rh001_022_002-    i_022    tia_h_in_001_002-    9434
Rh001_023_002+    i_023    tia_h_in_001_002+    15000
Rh001_023_002-    i_023    tia_h_in_001_002-    9238
Rh001_024_002+    i_024    tia_h_in_001_002+    15000
Rh001_024_002-    i_024    tia_h_in_001_002-    9216
Rh001_025_002+    i_025    tia_h_in_001_002+    15000
Rh001_025_002-    i_025    tia_h_in_001_002-    8930

* Neuron 3
Rh001_001_003+    i_001    tia_h_in_001_003+    15000
Rh001_001_003-    i_001    tia_h_in_001_003-    9425
Rh001_002_003+    i_002    tia_h_in_001_003+    15000
Rh001_002_003-    i_002    tia_h_in_001_003-    10070
Rh001_003_003+    i_003    tia_h_in_001_003+    15000
Rh001_003_003-    i_003    tia_h_in_001_003-    10130
Rh001_004_003+    i_004    tia_h_in_001_003+    15000
Rh001_004_003-    i_004    tia_h_in_001_003-    10130
Rh001_005_003+    i_005    tia_h_in_001_003+    15000
Rh001_005_003-    i_005    tia_h_in_001_003-    10221
Rh001_006_003+    i_006    tia_h_in_001_003+    15000
Rh001_006_003-    i_006    tia_h_in_001_003-    9853
Rh001_007_003+    i_007    tia_h_in_001_003+    15000
Rh001_007_003-    i_007    tia_h_in_001_003-    10038
Rh001_008_003+    i_008    tia_h_in_001_003+    15000
Rh001_008_003-    i_008    tia_h_in_001_003-    10175
Rh001_009_003+    i_009    tia_h_in_001_003+    15000
Rh001_009_003-    i_009    tia_h_in_001_003-    10304
Rh001_010_003+    i_010    tia_h_in_001_003+    15000
Rh001_010_003-    i_010    tia_h_in_001_003-    10291
Rh001_011_003+    i_011    tia_h_in_001_003+    15000
Rh001_011_003-    i_011    tia_h_in_001_003-    10506
Rh001_012_003+    i_012    tia_h_in_001_003+    15000
Rh001_012_003-    i_012    tia_h_in_001_003-    10234
Rh001_013_003+    i_013    tia_h_in_001_003+    15000
Rh001_013_003-    i_013    tia_h_in_001_003-    10558
Rh001_014_003+    i_014    tia_h_in_001_003+    15000
Rh001_014_003-    i_014    tia_h_in_001_003-    10156
Rh001_015_003+    i_015    tia_h_in_001_003+    15000
Rh001_015_003-    i_015    tia_h_in_001_003-    10194
Rh001_016_003+    i_016    tia_h_in_001_003+    15000
Rh001_016_003-    i_016    tia_h_in_001_003-    10311
Rh001_017_003+    i_017    tia_h_in_001_003+    15000
Rh001_017_003-    i_017    tia_h_in_001_003-    10608
Rh001_018_003+    i_018    tia_h_in_001_003+    15000
Rh001_018_003-    i_018    tia_h_in_001_003-    10280
Rh001_019_003+    i_019    tia_h_in_001_003+    15000
Rh001_019_003-    i_019    tia_h_in_001_003-    10236
Rh001_020_003+    i_020    tia_h_in_001_003+    15000
Rh001_020_003-    i_020    tia_h_in_001_003-    10059
Rh001_021_003+    i_021    tia_h_in_001_003+    15000
Rh001_021_003-    i_021    tia_h_in_001_003-    9911
Rh001_022_003+    i_022    tia_h_in_001_003+    15000
Rh001_022_003-    i_022    tia_h_in_001_003-    9952
Rh001_023_003+    i_023    tia_h_in_001_003+    15000
Rh001_023_003-    i_023    tia_h_in_001_003-    10227
Rh001_024_003+    i_024    tia_h_in_001_003+    15000
Rh001_024_003-    i_024    tia_h_in_001_003-    10168
Rh001_025_003+    i_025    tia_h_in_001_003+    15000
Rh001_025_003-    i_025    tia_h_in_001_003-    9709

* Neuron 4
Rh001_001_004+    i_001    tia_h_in_001_004+    13457
Rh001_001_004-    i_001    tia_h_in_001_004-    15000
Rh001_002_004+    i_002    tia_h_in_001_004+    15000
Rh001_002_004-    i_002    tia_h_in_001_004-    12997
Rh001_003_004+    i_003    tia_h_in_001_004+    15000
Rh001_003_004-    i_003    tia_h_in_001_004-    12632
Rh001_004_004+    i_004    tia_h_in_001_004+    14607
Rh001_004_004-    i_004    tia_h_in_001_004-    15000
Rh001_005_004+    i_005    tia_h_in_001_004+    15000
Rh001_005_004-    i_005    tia_h_in_001_004-    13271
Rh001_006_004+    i_006    tia_h_in_001_004+    13893
Rh001_006_004-    i_006    tia_h_in_001_004-    15000
Rh001_007_004+    i_007    tia_h_in_001_004+    15000
Rh001_007_004-    i_007    tia_h_in_001_004-    13958
Rh001_008_004+    i_008    tia_h_in_001_004+    14549
Rh001_008_004-    i_008    tia_h_in_001_004-    15000
Rh001_009_004+    i_009    tia_h_in_001_004+    15000
Rh001_009_004-    i_009    tia_h_in_001_004-    12174
Rh001_010_004+    i_010    tia_h_in_001_004+    15000
Rh001_010_004-    i_010    tia_h_in_001_004-    12874
Rh001_011_004+    i_011    tia_h_in_001_004+    15000
Rh001_011_004-    i_011    tia_h_in_001_004-    14527
Rh001_012_004+    i_012    tia_h_in_001_004+    14800
Rh001_012_004-    i_012    tia_h_in_001_004-    15000
Rh001_013_004+    i_013    tia_h_in_001_004+    15000
Rh001_013_004-    i_013    tia_h_in_001_004-    13328
Rh001_014_004+    i_014    tia_h_in_001_004+    13792
Rh001_014_004-    i_014    tia_h_in_001_004-    15000
Rh001_015_004+    i_015    tia_h_in_001_004+    13478
Rh001_015_004-    i_015    tia_h_in_001_004-    15000
Rh001_016_004+    i_016    tia_h_in_001_004+    15000
Rh001_016_004-    i_016    tia_h_in_001_004-    12571
Rh001_017_004+    i_017    tia_h_in_001_004+    15000
Rh001_017_004-    i_017    tia_h_in_001_004-    13070
Rh001_018_004+    i_018    tia_h_in_001_004+    13140
Rh001_018_004-    i_018    tia_h_in_001_004-    15000
Rh001_019_004+    i_019    tia_h_in_001_004+    15000
Rh001_019_004-    i_019    tia_h_in_001_004-    13434
Rh001_020_004+    i_020    tia_h_in_001_004+    15000
Rh001_020_004-    i_020    tia_h_in_001_004-    13561
Rh001_021_004+    i_021    tia_h_in_001_004+    15000
Rh001_021_004-    i_021    tia_h_in_001_004-    11906
Rh001_022_004+    i_022    tia_h_in_001_004+    15000
Rh001_022_004-    i_022    tia_h_in_001_004-    12878
Rh001_023_004+    i_023    tia_h_in_001_004+    15000
Rh001_023_004-    i_023    tia_h_in_001_004-    14969
Rh001_024_004+    i_024    tia_h_in_001_004+    15000
Rh001_024_004-    i_024    tia_h_in_001_004-    14183
Rh001_025_004+    i_025    tia_h_in_001_004+    15000
Rh001_025_004-    i_025    tia_h_in_001_004-    12559

* Neuron 5
Rh001_001_005+    i_001    tia_h_in_001_005+    15000
Rh001_001_005-    i_001    tia_h_in_001_005-    14856
Rh001_002_005+    i_002    tia_h_in_001_005+    9571
Rh001_002_005-    i_002    tia_h_in_001_005-    15000
Rh001_003_005+    i_003    tia_h_in_001_005+    9971
Rh001_003_005-    i_003    tia_h_in_001_005-    15000
Rh001_004_005+    i_004    tia_h_in_001_005+    9637
Rh001_004_005-    i_004    tia_h_in_001_005-    15000
Rh001_005_005+    i_005    tia_h_in_001_005+    9315
Rh001_005_005-    i_005    tia_h_in_001_005-    15000
Rh001_006_005+    i_006    tia_h_in_001_005+    10480
Rh001_006_005-    i_006    tia_h_in_001_005-    15000
Rh001_007_005+    i_007    tia_h_in_001_005+    7595
Rh001_007_005-    i_007    tia_h_in_001_005-    15000
Rh001_008_005+    i_008    tia_h_in_001_005+    8830
Rh001_008_005-    i_008    tia_h_in_001_005-    15000
Rh001_009_005+    i_009    tia_h_in_001_005+    8631
Rh001_009_005-    i_009    tia_h_in_001_005-    15000
Rh001_010_005+    i_010    tia_h_in_001_005+    9256
Rh001_010_005-    i_010    tia_h_in_001_005-    15000
Rh001_011_005+    i_011    tia_h_in_001_005+    7997
Rh001_011_005-    i_011    tia_h_in_001_005-    15000
Rh001_012_005+    i_012    tia_h_in_001_005+    9370
Rh001_012_005-    i_012    tia_h_in_001_005-    15000
Rh001_013_005+    i_013    tia_h_in_001_005+    9179
Rh001_013_005-    i_013    tia_h_in_001_005-    15000
Rh001_014_005+    i_014    tia_h_in_001_005+    9408
Rh001_014_005-    i_014    tia_h_in_001_005-    15000
Rh001_015_005+    i_015    tia_h_in_001_005+    7813
Rh001_015_005-    i_015    tia_h_in_001_005-    15000
Rh001_016_005+    i_016    tia_h_in_001_005+    8879
Rh001_016_005-    i_016    tia_h_in_001_005-    15000
Rh001_017_005+    i_017    tia_h_in_001_005+    8994
Rh001_017_005-    i_017    tia_h_in_001_005-    15000
Rh001_018_005+    i_018    tia_h_in_001_005+    9153
Rh001_018_005-    i_018    tia_h_in_001_005-    15000
Rh001_019_005+    i_019    tia_h_in_001_005+    8261
Rh001_019_005-    i_019    tia_h_in_001_005-    15000
Rh001_020_005+    i_020    tia_h_in_001_005+    10987
Rh001_020_005-    i_020    tia_h_in_001_005-    15000
Rh001_021_005+    i_021    tia_h_in_001_005+    9553
Rh001_021_005-    i_021    tia_h_in_001_005-    15000
Rh001_022_005+    i_022    tia_h_in_001_005+    9865
Rh001_022_005-    i_022    tia_h_in_001_005-    15000
Rh001_023_005+    i_023    tia_h_in_001_005+    9094
Rh001_023_005-    i_023    tia_h_in_001_005-    15000
Rh001_024_005+    i_024    tia_h_in_001_005+    9469
Rh001_024_005-    i_024    tia_h_in_001_005-    15000
Rh001_025_005+    i_025    tia_h_in_001_005+    13827
Rh001_025_005-    i_025    tia_h_in_001_005-    15000

* ----- Bias


Rb_h001_001+    b_001    tia_h_in_001_001+    8508
Rb_h001_001-    b_001    tia_h_in_001_001-    15000
Rb_h001_002+    b_001    tia_h_in_001_002+    5497
Rb_h001_002-    b_001    tia_h_in_001_002-    15000
Rb_h001_003+    b_001    tia_h_in_001_003+    6245
Rb_h001_003-    b_001    tia_h_in_001_003-    15000
Rb_h001_004+    b_001    tia_h_in_001_004+    15000
Rb_h001_004-    b_001    tia_h_in_001_004-    11427
Rb_h001_005+    b_001    tia_h_in_001_005+    15000
Rb_h001_005-    b_001    tia_h_in_001_005-    11053

* ----- Weights
* Layer 002

* Neuron 1
Rh002_001_001+    hidden_activ_out_h001_001    tia_h_in_002_001+    15000
Rh002_001_001-    hidden_activ_out_h001_001    tia_h_in_002_001-    8114
Rh002_002_001+    hidden_activ_out_h001_002    tia_h_in_002_001+    15000
Rh002_002_001-    hidden_activ_out_h001_002    tia_h_in_002_001-    5658
Rh002_003_001+    hidden_activ_out_h001_003    tia_h_in_002_001+    15000
Rh002_003_001-    hidden_activ_out_h001_003    tia_h_in_002_001-    5000
Rh002_004_001+    hidden_activ_out_h001_004    tia_h_in_002_001+    15000
Rh002_004_001-    hidden_activ_out_h001_004    tia_h_in_002_001-    9962
Rh002_005_001+    hidden_activ_out_h001_005    tia_h_in_002_001+    8147
Rh002_005_001-    hidden_activ_out_h001_005    tia_h_in_002_001-    15000

* ----- Bias


Rb_h002_001+    b_002    tia_h_in_002_001+    8887
Rb_h002_001-    b_002    tia_h_in_002_001-    15000


* ----- Difference (V(R+) - V(R-))

* Layer 000
* Neuron 1
Rh001_fb_001+     tia_h_in_001_001+ tia_h_out_001_001+ 4663.599371910095
Rh001_fb_001-     tia_h_in_001_001- tia_h_out_001_001- 4663.599371910095
XUh001_001+       0 tia_h_in_001_001+ Vcc+ Vcc- tia_h_out_001_001+ Ve OPA684_0
XUh001_001-       0 tia_h_in_001_001- Vcc+ Vcc- tia_h_out_001_001- Ve OPA684_0
Rh001_sum_001+    tia_h_out_001_001+ sum_h_in_001_001- 260
Rh001_sum_001-    tia_h_out_001_001- sum_h_in_001_001+ 260
Rh001_sum_l_001   sum_h_in_001_001+ 0 650.0
Rh001_sum_fb_001  sum_h_in_001_001- sum_h_out_001_001 650.0
XUh001_sum_001    sum_h_in_001_001+ sum_h_in_001_001- Vcc+ Vcc- sum_h_out_001_001 MAX4223
* Neuron 2
Rh001_fb_002+     tia_h_in_001_002+ tia_h_out_001_002+ 4663.599371910095
Rh001_fb_002-     tia_h_in_001_002- tia_h_out_001_002- 4663.599371910095
XUh001_002+       0 tia_h_in_001_002+ Vcc+ Vcc- tia_h_out_001_002+ Ve OPA684_0
XUh001_002-       0 tia_h_in_001_002- Vcc+ Vcc- tia_h_out_001_002- Ve OPA684_0
Rh001_sum_002+    tia_h_out_001_002+ sum_h_in_001_002- 260
Rh001_sum_002-    tia_h_out_001_002- sum_h_in_001_002+ 260
Rh001_sum_l_002   sum_h_in_001_002+ 0 650.0
Rh001_sum_fb_002  sum_h_in_001_002- sum_h_out_001_002 650.0
XUh001_sum_002    sum_h_in_001_002+ sum_h_in_001_002- Vcc+ Vcc- sum_h_out_001_002 MAX4223
* Neuron 3
Rh001_fb_003+     tia_h_in_001_003+ tia_h_out_001_003+ 4663.599371910095
Rh001_fb_003-     tia_h_in_001_003- tia_h_out_001_003- 4663.599371910095
XUh001_003+       0 tia_h_in_001_003+ Vcc+ Vcc- tia_h_out_001_003+ Ve OPA684_0
XUh001_003-       0 tia_h_in_001_003- Vcc+ Vcc- tia_h_out_001_003- Ve OPA684_0
Rh001_sum_003+    tia_h_out_001_003+ sum_h_in_001_003- 260
Rh001_sum_003-    tia_h_out_001_003- sum_h_in_001_003+ 260
Rh001_sum_l_003   sum_h_in_001_003+ 0 650.0
Rh001_sum_fb_003  sum_h_in_001_003- sum_h_out_001_003 650.0
XUh001_sum_003    sum_h_in_001_003+ sum_h_in_001_003- Vcc+ Vcc- sum_h_out_001_003 MAX4223
* Neuron 4
Rh001_fb_004+     tia_h_in_001_004+ tia_h_out_001_004+ 4663.599371910095
Rh001_fb_004-     tia_h_in_001_004- tia_h_out_001_004- 4663.599371910095
XUh001_004+       0 tia_h_in_001_004+ Vcc+ Vcc- tia_h_out_001_004+ Ve OPA684_0
XUh001_004-       0 tia_h_in_001_004- Vcc+ Vcc- tia_h_out_001_004- Ve OPA684_0
Rh001_sum_004+    tia_h_out_001_004+ sum_h_in_001_004- 260
Rh001_sum_004-    tia_h_out_001_004- sum_h_in_001_004+ 260
Rh001_sum_l_004   sum_h_in_001_004+ 0 650.0
Rh001_sum_fb_004  sum_h_in_001_004- sum_h_out_001_004 650.0
XUh001_sum_004    sum_h_in_001_004+ sum_h_in_001_004- Vcc+ Vcc- sum_h_out_001_004 MAX4223
* Neuron 5
Rh001_fb_005+     tia_h_in_001_005+ tia_h_out_001_005+ 4663.599371910095
Rh001_fb_005-     tia_h_in_001_005- tia_h_out_001_005- 4663.599371910095
XUh001_005+       0 tia_h_in_001_005+ Vcc+ Vcc- tia_h_out_001_005+ Ve OPA684_0
XUh001_005-       0 tia_h_in_001_005- Vcc+ Vcc- tia_h_out_001_005- Ve OPA684_0
Rh001_sum_005+    tia_h_out_001_005+ sum_h_in_001_005- 260
Rh001_sum_005-    tia_h_out_001_005- sum_h_in_001_005+ 260
Rh001_sum_l_005   sum_h_in_001_005+ 0 650.0
Rh001_sum_fb_005  sum_h_in_001_005- sum_h_out_001_005 650.0
XUh001_sum_005    sum_h_in_001_005+ sum_h_in_001_005- Vcc+ Vcc- sum_h_out_001_005 MAX4223

* Layer 001
* Neuron 1
Rh002_fb_001+     tia_h_in_002_001+ tia_h_out_002_001+ 4663.599371910095
Rh002_fb_001-     tia_h_in_002_001- tia_h_out_002_001- 4663.599371910095
XUh002_001+       0 tia_h_in_002_001+ Vcc+ Vcc- tia_h_out_002_001+ Ve OPA684_0
XUh002_001-       0 tia_h_in_002_001- Vcc+ Vcc- tia_h_out_002_001- Ve OPA684_0
Rh002_sum_001+    tia_h_out_002_001+ sum_h_in_002_001- 260
Rh002_sum_001-    tia_h_out_002_001- sum_h_in_002_001+ 260
Rh002_sum_l_001   sum_h_in_002_001+ 0 650.0
Rh002_sum_fb_001  sum_h_in_002_001- sum_h_out_002_001 650.0
XUh002_sum_001    sum_h_in_002_001+ sum_h_in_002_001- Vcc+ Vcc- sum_h_out_002_001 MAX4223


* ----- Activation function Hard-Tanh)


* Layer 000
* Neuron 1
* XHardTanh_h001_001 sum_h_out_001_001 hidden_activ_out_h001_001 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_001 sum_h_out_001_001 hidden_activ_out_h001_001 ReLU
* Neuron 2
* XHardTanh_h001_002 sum_h_out_001_002 hidden_activ_out_h001_002 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_002 sum_h_out_001_002 hidden_activ_out_h001_002 ReLU
* Neuron 3
* XHardTanh_h001_003 sum_h_out_001_003 hidden_activ_out_h001_003 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_003 sum_h_out_001_003 hidden_activ_out_h001_003 ReLU
* Neuron 4
* XHardTanh_h001_004 sum_h_out_001_004 hidden_activ_out_h001_004 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_004 sum_h_out_001_004 hidden_activ_out_h001_004 ReLU
* Neuron 5
* XHardTanh_h001_005 sum_h_out_001_005 hidden_activ_out_h001_005 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_001_005 sum_h_out_001_005 hidden_activ_out_h001_005 ReLU

* Layer 001
* Neuron 1
* XHardTanh_h002_001 sum_h_out_002_001 hidden_activ_out_h002_001 HardTanh PARAMS: V_clip=-0.39999999999999997
XReLU_002_001 sum_h_out_002_001 hidden_activ_out_h002_001 ReLU


.END
